*GAP co-working with Royal Road test chip simulation  

*Options
*.param hsimveriloga="RAM.va"
*.param hsimveriloga="RoyalRoad.va"
.hdl "RAM.va"
.hdl "RoyalRoad.va"
*.param hsimvdd=1.8
*.param hsimspeed=3
*.param hsimanalog=1.5
.probe v(*)	level=2	***** tran
.probe I(vdd)		***** tran

***CustomSim Parameters
.option XA_CMD="set_sim_level -level	6"
.option XA_CMD="set_save_state  -period_wall_time	12"

.lib	'hm1816m020233v11.lib'	tt	

.tran	20p	16u	*UIC	*sweep monte=30
*.option post		*post_version=2001	posttop=3	*list=element	*modmonte=1
*.option runlvl=1
*.option converge=5
*.store	repeat=7200

*Sources
vdd	vdd	0	1.8
.global	vdd

vMaster-Slave-Select-Pin-1-1	Master-Slave-Select-Pin-1-1	0	0	*Master
vMaster-Slave-Select-Pin-0-1	Master-Slave-Select-Pin-0-1	0	1.8

vMaster-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-1-2	0	1.8	*Slave
vMaster-Slave-Select-Pin-0-2	Master-Slave-Select-Pin-0-2	0	0

vMaster-Slave-Select-Pin-1-3	Master-Slave-Select-Pin-1-3	0	1.8	*Last Slave
vMaster-Slave-Select-Pin-0-3	Master-Slave-Select-Pin-0-3	0	1.8

vChromosome-Resolution-Pin	Chromosome-Resolution-Pin	0	1.8	*32 bits
vFitness-Resolution-Pin	Fitness-Resolution-Pin	0	0	*16 bits

vBest-Found-Emmigration-Pin	Best-Found-Emmigration-Pin	0	0	*First Offspring Sending

vNo-Elitism-Pin	No-Elitism-Pin	0	0	*Elitism Enabled

vDual-Ram-Pin	Dual-Ram-Pin	0	0	*Dual-Population Enabled

vRestart-Pin	Restart-Pin	0	pulse(0	1.8	0n	50p	50p	1n	100u)	*Restart at First Only
vStop-Pin	Stop-Pin	0	0	*No Stop in Process

vClock-1-Pin	Clock-1-Pin	0	pulse(0	1.8	0n	50p	50p	1.05n	2.2n)	*Main Clock
vClock-2-Pin	Clock-2-Pin	0	pulse(0	1.8	0n	50p	50p	0.6n	1.3n)	*Second Clock for Parallel Processing

vPopulation-Size-Pin-0	Population-Size-Pin-0	0	1.8	*256
vPopulation-Size-Pin-1	Population-Size-Pin-1	0	1.8

vRandom-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-1	0	1.8	*Every 2 Iterations
vRandom-Immigrants-Gap-Pin-0	Random-Immigrants-Gap-Pin-0	0	0

vMutation-Rate-Pin-0	Mutation-Rate-Pin-0	0	0
vMutation-Rate-Pin-1	Mutation-Rate-Pin-1	0	1.8
vMutation-Rate-Pin-2	Mutation-Rate-Pin-2	0	0
vMutation-Rate-Pin-3	Mutation-Rate-Pin-3	0	1.8
vMutation-Rate-Pin-4	Mutation-Rate-Pin-4	0	0	*11/128
vMutation-Rate-Pin-5	Mutation-Rate-Pin-5	0	0
vMutation-Rate-Pin-6	Mutation-Rate-Pin-6	0	0

vCrossover-Rate-Pin-0	Crossover-Rate-Pin-0	0	0
vCrossover-Rate-Pin-1	Crossover-Rate-Pin-1	0	0
vCrossover-Rate-Pin-2	Crossover-Rate-Pin-2	0	0	*89/128
vCrossover-Rate-Pin-3	Crossover-Rate-Pin-3	0	1.8
vCrossover-Rate-Pin-4	Crossover-Rate-Pin-4	0	1.8
vCrossover-Rate-Pin-5	Crossover-Rate-Pin-5	0	0
vCrossover-Rate-Pin-6	Crossover-Rate-Pin-6	0	1.8

vMigration-Gap-Pin-1	Migration-Gap-Pin-1	0	1.8	*Every 4 Iterations
vMigration-Gap-Pin-0	Migration-Gap-Pin-0	0	1.8

vSecond-SPI-Ready-Pin	Second-SPI-Ready-Pin	0	1.8	*Second Immigration Module is Active

vFitness-or-Cost-Pin	Fitness-or-Cost-Pin	0	1.8	*Cost

vTournament-Size-Pin-1	Tournament-Size-Pin-1	0	1.8
vTournament-Size-Pin-0	Tournament-Size-Pin-0	0	1.8	*16

vIteration-Number-Pin-0	Iteration-Number-Pin-0	0	0
vIteration-Number-Pin-1	Iteration-Number-Pin-1	0	0	*256
vIteration-Number-Pin-2	Iteration-Number-Pin-2	0	1.8

vUniform-Mutation-Pin	Uniform-Mutation-Pin	0	1.8	*Uniform Mutation
vOne-Point-Mutation-Pin	One-Point-Mutation-Pin	0	0

vUniform-Crossover-Pin	Uniform-Crossover-Pin	0	1.8	*Uniform Crossover
vCrossover-Type-Pin-1	Crossover-Type-Pin-1	0	0
vCrossover-Type-Pin-0	Crossover-Type-Pin-0	0	0

vPipeline-Stages-Pin-3	Pipeline-Stages-Pin-3	0	0
vPipeline-Stages-Pin-2	Pipeline-Stages-Pin-2	0	1.8
vPipeline-Stages-Pin-1	Pipeline-Stages-Pin-1	0	0	*Five Pipeline Stages Latency in TWO FU STRUCTURE
vPipeline-Stages-Pin-0	Pipeline-Stages-Pin-0	0	1.8

vCrossover-In-Req-Pin	Crossover-In-Req-Pin	0	0	*No Crossover State Transmission in Uniform Crossover
vCrossover-In-Data-Pin	Crossover-In-Data-Pin	0	0
vCrossover-Out-Ack-Pin	Crossover-Out-Ack-Pin	0	0

*vSPI-In1-Line1	SPI-In1-Line1	0	0
*vSPI-In1-Line2	SPI-In1-Line2	0	0
*vSPI-In1-Line3	SPI-In1-Line3	0	0
*vSPI-In1-Line4	SPI-In1-Line4	0	0
*vSPI-In1-clk-Pin	SPI-In1-clk-Pin	0	0
*vSPI-In1-CS-Pin	SPI-In1-CS-Pin	0	0

*vSPI-In2-Line1	SPI-In2-Line1	0	0
*vSPI-In2-Line2	SPI-In2-Line2	0	0
*vSPI-In2-Line3	SPI-In2-Line3	0	0
*vSPI-In2-Line4	SPI-In2-Line4	0	0
*vSPI-In2-clk-Pin	SPI-In2-clk-Pin	0	0
*vSPI-In2-CS-Pin	SPI-In2-CS-Pin	0	0

vFitness-Estimation-Discard-Pin	Fitness-Estimation-Discard-Pin	0	0	*No Discard Operator

vPRNG-Seed-Select-Pin-0-1	PRNG-Seed-Select-Pin-0-1	0	0	*1st PRNG Seed
vPRNG-Seed-Select-Pin-1-1	PRNG-Seed-Select-Pin-1-1	0	0
vPRNG-Seed-Select-Pin-2-1	PRNG-Seed-Select-Pin-2-1	0	0
vPRNG-Seed-Select-Pin-3-1	PRNG-Seed-Select-Pin-3-1	0	0

vPRNG-Seed-Select-Pin-0-2	PRNG-Seed-Select-Pin-0-2	0	1.8	*2nd PRNG Seed
vPRNG-Seed-Select-Pin-1-2	PRNG-Seed-Select-Pin-1-2	0	0
vPRNG-Seed-Select-Pin-2-2	PRNG-Seed-Select-Pin-2-2	0	0
vPRNG-Seed-Select-Pin-3-2	PRNG-Seed-Select-Pin-3-2	0	0

vPRNG-Seed-Select-Pin-0-3	PRNG-Seed-Select-Pin-0-3	0	0	*3rd PRNG Seed
vPRNG-Seed-Select-Pin-1-3	PRNG-Seed-Select-Pin-1-3	0	1.8
vPRNG-Seed-Select-Pin-2-3	PRNG-Seed-Select-Pin-2-3	0	0
vPRNG-Seed-Select-Pin-3-3	PRNG-Seed-Select-Pin-3-3	0	0

vPRNG-Seed-Select-Pin-0-4	PRNG-Seed-Select-Pin-0-4	0	1.8	*4th PRNG Seed
vPRNG-Seed-Select-Pin-1-4	PRNG-Seed-Select-Pin-1-4	0	1.8
vPRNG-Seed-Select-Pin-2-4	PRNG-Seed-Select-Pin-2-4	0	0
vPRNG-Seed-Select-Pin-3-4	PRNG-Seed-Select-Pin-3-4	0	0

vPRNG-Seed-Select-Pin-0-5	PRNG-Seed-Select-Pin-0-5	0	0	*5th PRNG Seed
vPRNG-Seed-Select-Pin-1-5	PRNG-Seed-Select-Pin-1-5	0	0
vPRNG-Seed-Select-Pin-2-5	PRNG-Seed-Select-Pin-2-5	0	1.8
vPRNG-Seed-Select-Pin-3-5	PRNG-Seed-Select-Pin-3-5	0	0

vPRNG-Seed-Select-Pin-0-6	PRNG-Seed-Select-Pin-0-6	0	1.8	*6th PRNG Seed
vPRNG-Seed-Select-Pin-1-6	PRNG-Seed-Select-Pin-1-6	0	0
vPRNG-Seed-Select-Pin-2-6	PRNG-Seed-Select-Pin-2-6	0	1.8
vPRNG-Seed-Select-Pin-3-6	PRNG-Seed-Select-Pin-3-6	0	0

vPRNG-Seed-Select-Pin-0-7	PRNG-Seed-Select-Pin-0-7	0	0	*7th PRNG Seed
vPRNG-Seed-Select-Pin-1-7	PRNG-Seed-Select-Pin-1-7	0	1.8
vPRNG-Seed-Select-Pin-2-7	PRNG-Seed-Select-Pin-2-7	0	1.8
vPRNG-Seed-Select-Pin-3-7	PRNG-Seed-Select-Pin-3-7	0	0

vPRNG-Seed-Select-Pin-0-8	PRNG-Seed-Select-Pin-0-8	0	1.8	*8th PRNG Seed
vPRNG-Seed-Select-Pin-1-8	PRNG-Seed-Select-Pin-1-8	0	1.8
vPRNG-Seed-Select-Pin-2-8	PRNG-Seed-Select-Pin-2-8	0	1.8
vPRNG-Seed-Select-Pin-3-8	PRNG-Seed-Select-Pin-3-8	0	0

vPRNG-Seed-Select-Pin-0-9	PRNG-Seed-Select-Pin-0-9	0	0	*9th PRNG Seed
vPRNG-Seed-Select-Pin-1-9	PRNG-Seed-Select-Pin-1-9	0	0
vPRNG-Seed-Select-Pin-2-9	PRNG-Seed-Select-Pin-2-9	0	0
vPRNG-Seed-Select-Pin-3-9	PRNG-Seed-Select-Pin-3-9	0	1.8

vPRNG-Seed-Select-Pin-0-10	PRNG-Seed-Select-Pin-0-10	0	1.8	*10th PRNG Seed
vPRNG-Seed-Select-Pin-1-10	PRNG-Seed-Select-Pin-1-10	0	0
vPRNG-Seed-Select-Pin-2-10	PRNG-Seed-Select-Pin-2-10	0	0
vPRNG-Seed-Select-Pin-3-10	PRNG-Seed-Select-Pin-3-10	0	1.8

vPRNG-Seed-Select-Pin-0-11	PRNG-Seed-Select-Pin-0-11	0	0	*11th PRNG Seed
vPRNG-Seed-Select-Pin-1-11	PRNG-Seed-Select-Pin-1-11	0	1.8
vPRNG-Seed-Select-Pin-2-11	PRNG-Seed-Select-Pin-2-11	0	0
vPRNG-Seed-Select-Pin-3-11	PRNG-Seed-Select-Pin-3-11	0	1.8

vPRNG-Seed-Select-Pin-0-12	PRNG-Seed-Select-Pin-0-12	0	1.8	*12th PRNG Seed
vPRNG-Seed-Select-Pin-1-12	PRNG-Seed-Select-Pin-1-12	0	1.8
vPRNG-Seed-Select-Pin-2-12	PRNG-Seed-Select-Pin-2-12	0	0
vPRNG-Seed-Select-Pin-3-12	PRNG-Seed-Select-Pin-3-12	0	1.8

vPRNG-Seed-Select-Pin-0-13	PRNG-Seed-Select-Pin-0-13	0	0	*13th PRNG Seed
vPRNG-Seed-Select-Pin-1-13	PRNG-Seed-Select-Pin-1-13	0	0
vPRNG-Seed-Select-Pin-2-13	PRNG-Seed-Select-Pin-2-13	0	1.8
vPRNG-Seed-Select-Pin-3-13	PRNG-Seed-Select-Pin-3-13	0	1.8

vPRNG-Seed-Select-Pin-0-14	PRNG-Seed-Select-Pin-0-14	0	1.8	*14th PRNG Seed
vPRNG-Seed-Select-Pin-1-14	PRNG-Seed-Select-Pin-1-14	0	0
vPRNG-Seed-Select-Pin-2-14	PRNG-Seed-Select-Pin-2-14	0	1.8
vPRNG-Seed-Select-Pin-3-14	PRNG-Seed-Select-Pin-3-14	0	1.8

vPRNG-Seed-Select-Pin-0-15	PRNG-Seed-Select-Pin-0-15	0	0	*15th PRNG Seed
vPRNG-Seed-Select-Pin-1-15	PRNG-Seed-Select-Pin-1-15	0	1.8
vPRNG-Seed-Select-Pin-2-15	PRNG-Seed-Select-Pin-2-15	0	1.8
vPRNG-Seed-Select-Pin-3-15	PRNG-Seed-Select-Pin-3-15	0	1.8

vPRNG-Seed-Select-Pin-0-16	PRNG-Seed-Select-Pin-0-16	0	1.8	*16th PRNG Seed
vPRNG-Seed-Select-Pin-1-16	PRNG-Seed-Select-Pin-1-16	0	1.8
vPRNG-Seed-Select-Pin-2-16	PRNG-Seed-Select-Pin-2-16	0	1.8
vPRNG-Seed-Select-Pin-3-16	PRNG-Seed-Select-Pin-3-16	0	1.8


*GAPs
*names are based on the master chip namings
x1	Master-Slave-Select-Pin-1-1	Master-Slave-Select-Pin-0-1	Selection-Req-Pad1	Selection-Ack-Pin1-1	Address-Port-1-1	Address-Port-2-1	Address-Port-3-1	Address-Port-4-1	Address-Port-5-1	Address-Port-6-1	Address-Port-7-1	Address-Port-8-1	Address-Port-9-Elite-Selected-1	RNG-Pad-0-1-1	RNG-Pad-1-1-1	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-1-1	Crossover-Out-Data-Pad-1-1	Crossover-In-Ack-Pad-1-1	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-1-1	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad1-1	SPI-Out-Line2-Pad1-1	SPI-Out-Line3-Pad1-1	SPI-Out-Line4-Pad1-1	SPI-Out-clk-Pad1-1	SPI-Out-CS-Pad1-1	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad1-4	SPI-Out-Line2-Pad1-4	SPI-Out-Line3-Pad1-4	SPI-Out-Line4-Pad1-4	SPI-Out-clk-Pad1-4	SPI-Out-CS-Pad1-4	SPI-Out-Line1-Pad1-2	SPI-Out-Line2-Pad1-2	SPI-Out-Line3-Pad1-2	SPI-Out-Line4-Pad1-2	SPI-Out-clk-Pad1-2	SPI-Out-CS-Pad1-2	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-1	PRNG-Seed-Select-Pin-1-1	PRNG-Seed-Select-Pin-2-1	PRNG-Seed-Select-Pin-3-1	Fitness-Estimation-Ack-Pin-1	Fitness-Estimation-Req1-Pad1-1	Fitness-Estimation-Req2-Pad1-1	Fitness-Estimation-Ready1-Pad1-1	Fitness-Estimation-Ready2-Pad1-1	Fitness-Estimation-Discard-Pin	Data0-1	Data1-1	Data2-1	Data3-1	Data4-1	Data5-1	Data6-1	Data7-1	Data8-1	Data9-1	Data10-1	Data11-1	Data12-1	Data13-1	Data14-1	Data15-1	Data16-1	Data17-1	Data18-1	Data19-1	Data20-1	Data21-1	Data22-1	Data23-1	Data24-1	Data25-1	Data26-1	Data27-1	Data28-1	Data29-1	Data30-1	Data31-1	GAP
x2	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin2-1	Selection-Req-Pad1	Address-Port-1-1	Address-Port-2-1	Address-Port-3-1	Address-Port-4-1	Address-Port-5-1	Address-Port-6-1	Address-Port-7-1	Address-Port-8-1	Address-Port-9-Elite-Selected-1	RNG-Pad-0-2-1	RNG-Pad-1-2-1	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-2-1	Crossover-Out-Data-Pad-2-1	Crossover-In-Ack-Pad-2-1	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-2-1	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad2-1	SPI-Out-Line2-Pad2-1	SPI-Out-Line3-Pad2-1	SPI-Out-Line4-Pad2-1	SPI-Out-clk-Pad2-1	SPI-Out-CS-Pad2-1	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad2-4	SPI-Out-Line2-Pad2-4	SPI-Out-Line3-Pad2-4	SPI-Out-Line4-Pad2-4	SPI-Out-clk-Pad2-4	SPI-Out-CS-Pad2-4	SPI-Out-Line1-Pad2-2	SPI-Out-Line2-Pad2-2	SPI-Out-Line3-Pad2-2	SPI-Out-Line4-Pad2-2	SPI-Out-clk-Pad2-2	SPI-Out-CS-Pad2-2	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-2	PRNG-Seed-Select-Pin-1-2	PRNG-Seed-Select-Pin-2-2	PRNG-Seed-Select-Pin-3-2	Fitness-Estimation-Ack-Pin-1	Fitness-Estimation-Req1-Pad2-1	Fitness-Estimation-Req2-Pad2-1	Fitness-Estimation-Ready1-Pad2-1	Fitness-Estimation-Ready2-Pad2-1	Fitness-Estimation-Discard-Pin	Data32-1	Data33-1	Data34-1	Data35-1	Data36-1	Data37-1	Data38-1	Data39-1	Data40-1	Data41-1	Data42-1	Data43-1	Data44-1	Data45-1	Data46-1	Data47-1	Data48-1	Data49-1	Data50-1	Data51-1	Data52-1	Data53-1	Data54-1	Data55-1	Data56-1	Data57-1	Data58-1	Data59-1	Data60-1	Data61-1	Data62-1	Data63-1	GAP
x3	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin3-1	Selection-Req-Pad1	Address-Port-1-1	Address-Port-2-1	Address-Port-3-1	Address-Port-4-1	Address-Port-5-1	Address-Port-6-1	Address-Port-7-1	Address-Port-8-1	Address-Port-9-Elite-Selected-1	RNG-Pad-0-3-1	RNG-Pad-1-3-1	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-3-1	Crossover-Out-Data-Pad-3-1	Crossover-In-Ack-Pad-3-1	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-3-1	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad3-1	SPI-Out-Line2-Pad3-1	SPI-Out-Line3-Pad3-1	SPI-Out-Line4-Pad3-1	SPI-Out-clk-Pad3-1	SPI-Out-CS-Pad3-1	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad3-4	SPI-Out-Line2-Pad3-4	SPI-Out-Line3-Pad3-4	SPI-Out-Line4-Pad3-4	SPI-Out-clk-Pad3-4	SPI-Out-CS-Pad3-4	SPI-Out-Line1-Pad3-2	SPI-Out-Line2-Pad3-2	SPI-Out-Line3-Pad3-2	SPI-Out-Line4-Pad3-2	SPI-Out-clk-Pad3-2	SPI-Out-CS-Pad3-2	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-3	PRNG-Seed-Select-Pin-1-3	PRNG-Seed-Select-Pin-2-3	PRNG-Seed-Select-Pin-3-3	Fitness-Estimation-Ack-Pin-1	Fitness-Estimation-Req1-Pad3-1	Fitness-Estimation-Req2-Pad3-1	Fitness-Estimation-Ready1-Pad3-1	Fitness-Estimation-Ready2-Pad3-1	Fitness-Estimation-Discard-Pin	Data64-1	Data65-1	Data66-1	Data67-1	Data68-1	Data69-1	Data70-1	Data71-1	Data72-1	Data73-1	Data74-1	Data75-1	Data76-1	Data77-1	Data78-1	Data79-1	Data80-1	Data81-1	Data82-1	Data83-1	Data84-1	Data85-1	Data86-1	Data87-1	Data88-1	Data89-1	Data90-1	Data91-1	Data92-1	Data93-1	Data94-1	Data95-1	GAP
x4	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin4-1	Selection-Req-Pad1	Address-Port-1-1	Address-Port-2-1	Address-Port-3-1	Address-Port-4-1	Address-Port-5-1	Address-Port-6-1	Address-Port-7-1	Address-Port-8-1	Address-Port-9-Elite-Selected-1	RNG-Pad-0-4-1	RNG-Pad-1-4-1	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-4-1	Crossover-Out-Data-Pad-4-1	Crossover-In-Ack-Pad-4-1	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-4-1	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad4-1	SPI-Out-Line2-Pad4-1	SPI-Out-Line3-Pad4-1	SPI-Out-Line4-Pad4-1	SPI-Out-clk-Pad4-1	SPI-Out-CS-Pad4-1	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad4-4	SPI-Out-Line2-Pad4-4	SPI-Out-Line3-Pad4-4	SPI-Out-Line4-Pad4-4	SPI-Out-clk-Pad4-4	SPI-Out-CS-Pad4-4	SPI-Out-Line1-Pad4-2	SPI-Out-Line2-Pad4-2	SPI-Out-Line3-Pad4-2	SPI-Out-Line4-Pad4-2	SPI-Out-clk-Pad4-2	SPI-Out-CS-Pad4-2	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-4	PRNG-Seed-Select-Pin-1-4	PRNG-Seed-Select-Pin-2-4	PRNG-Seed-Select-Pin-3-4	Fitness-Estimation-Ack-Pin-1	Fitness-Estimation-Req1-Pad4-1	Fitness-Estimation-Req2-Pad4-1	Fitness-Estimation-Ready1-Pad4-1	Fitness-Estimation-Ready2-Pad4-1	Fitness-Estimation-Discard-Pin	Data96-1	Data97-1	Data98-1	Data99-1	Data100-1	Data101-1	Data102-1	Data103-1	Data104-1	Data105-1	Data106-1	Data107-1	Data108-1	Data109-1	Data110-1	Data111-1	Data112-1	Data113-1	Data114-1	Data115-1	Data116-1	Data117-1	Data118-1	Data119-1	Data120-1	Data121-1	Data122-1	Data123-1	Data124-1	Data125-1	Data126-1	Data127-1	GAP
x5	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin5-1	Selection-Req-Pad1	Address-Port-1-1	Address-Port-2-1	Address-Port-3-1	Address-Port-4-1	Address-Port-5-1	Address-Port-6-1	Address-Port-7-1	Address-Port-8-1	Address-Port-9-Elite-Selected-1	RNG-Pad-0-5-1	RNG-Pad-1-5-1	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-5-1	Crossover-Out-Data-Pad-5-1	Crossover-In-Ack-Pad-5-1	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-5-1	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad5-1	SPI-Out-Line2-Pad5-1	SPI-Out-Line3-Pad5-1	SPI-Out-Line4-Pad5-1	SPI-Out-clk-Pad5-1	SPI-Out-CS-Pad5-1	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad5-4	SPI-Out-Line2-Pad5-4	SPI-Out-Line3-Pad5-4	SPI-Out-Line4-Pad5-4	SPI-Out-clk-Pad5-4	SPI-Out-CS-Pad5-4	SPI-Out-Line1-Pad5-2	SPI-Out-Line2-Pad5-2	SPI-Out-Line3-Pad5-2	SPI-Out-Line4-Pad5-2	SPI-Out-clk-Pad5-2	SPI-Out-CS-Pad5-2	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-5	PRNG-Seed-Select-Pin-1-5	PRNG-Seed-Select-Pin-2-5	PRNG-Seed-Select-Pin-3-5	Fitness-Estimation-Ack-Pin-1	Fitness-Estimation-Req1-Pad5-1	Fitness-Estimation-Req2-Pad5-1	Fitness-Estimation-Ready1-Pad5-1	Fitness-Estimation-Ready2-Pad5-1	Fitness-Estimation-Discard-Pin	Data128-1	Data129-1	Data130-1	Data131-1	Data132-1	Data133-1	Data134-1	Data135-1	Data136-1	Data137-1	Data138-1	Data139-1	Data140-1	Data141-1	Data142-1	Data143-1	Data144-1	Data145-1	Data146-1	Data147-1	Data148-1	Data149-1	Data150-1	Data151-1	Data152-1	Data153-1	Data154-1	Data155-1	Data156-1	Data157-1	Data158-1	Data159-1	GAP
x6	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin6-1	Selection-Req-Pad1	Address-Port-1-1	Address-Port-2-1	Address-Port-3-1	Address-Port-4-1	Address-Port-5-1	Address-Port-6-1	Address-Port-7-1	Address-Port-8-1	Address-Port-9-Elite-Selected-1	RNG-Pad-0-6-1	RNG-Pad-1-6-1	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-6-1	Crossover-Out-Data-Pad-6-1	Crossover-In-Ack-Pad-6-1	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-6-1	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad6-1	SPI-Out-Line2-Pad6-1	SPI-Out-Line3-Pad6-1	SPI-Out-Line4-Pad6-1	SPI-Out-clk-Pad6-1	SPI-Out-CS-Pad6-1	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad6-4	SPI-Out-Line2-Pad6-4	SPI-Out-Line3-Pad6-4	SPI-Out-Line4-Pad6-4	SPI-Out-clk-Pad6-4	SPI-Out-CS-Pad6-4	SPI-Out-Line1-Pad6-2	SPI-Out-Line2-Pad6-2	SPI-Out-Line3-Pad6-2	SPI-Out-Line4-Pad6-2	SPI-Out-clk-Pad6-2	SPI-Out-CS-Pad6-2	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-6	PRNG-Seed-Select-Pin-1-6	PRNG-Seed-Select-Pin-2-6	PRNG-Seed-Select-Pin-3-6	Fitness-Estimation-Ack-Pin-1	Fitness-Estimation-Req1-Pad6-1	Fitness-Estimation-Req2-Pad6-1	Fitness-Estimation-Ready1-Pad6-1	Fitness-Estimation-Ready2-Pad6-1	Fitness-Estimation-Discard-Pin	Data160-1	Data161-1	Data162-1	Data163-1	Data164-1	Data165-1	Data166-1	Data167-1	Data168-1	Data169-1	Data170-1	Data171-1	Data172-1	Data173-1	Data174-1	Data175-1	Data176-1	Data177-1	Data178-1	Data179-1	Data180-1	Data181-1	Data182-1	Data183-1	Data184-1	Data185-1	Data186-1	Data187-1	Data188-1	Data189-1	Data190-1	Data191-1	GAP
x7	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin7-1	Selection-Req-Pad1	Address-Port-1-1	Address-Port-2-1	Address-Port-3-1	Address-Port-4-1	Address-Port-5-1	Address-Port-6-1	Address-Port-7-1	Address-Port-8-1	Address-Port-9-Elite-Selected-1	RNG-Pad-0-7-1	RNG-Pad-1-7-1	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-7-1	Crossover-Out-Data-Pad-7-1	Crossover-In-Ack-Pad-7-1	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-7-1	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad7-1	SPI-Out-Line2-Pad7-1	SPI-Out-Line3-Pad7-1	SPI-Out-Line4-Pad7-1	SPI-Out-clk-Pad7-1	SPI-Out-CS-Pad7-1	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad7-4	SPI-Out-Line2-Pad7-4	SPI-Out-Line3-Pad7-4	SPI-Out-Line4-Pad7-4	SPI-Out-clk-Pad7-4	SPI-Out-CS-Pad7-4	SPI-Out-Line1-Pad7-2	SPI-Out-Line2-Pad7-2	SPI-Out-Line3-Pad7-2	SPI-Out-Line4-Pad7-2	SPI-Out-clk-Pad7-2	SPI-Out-CS-Pad7-2	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-7	PRNG-Seed-Select-Pin-1-7	PRNG-Seed-Select-Pin-2-7	PRNG-Seed-Select-Pin-3-7	Fitness-Estimation-Ack-Pin-1	Fitness-Estimation-Req1-Pad7-1	Fitness-Estimation-Req2-Pad7-1	Fitness-Estimation-Ready1-Pad7-1	Fitness-Estimation-Ready2-Pad7-1	Fitness-Estimation-Discard-Pin	Data192-1	Data193-1	Data194-1	Data195-1	Data196-1	Data197-1	Data198-1	Data199-1	Data200-1	Data201-1	Data202-1	Data203-1	Data204-1	Data205-1	Data206-1	Data207-1	Data208-1	Data209-1	Data210-1	Data211-1	Data212-1	Data213-1	Data214-1	Data215-1	Data216-1	Data217-1	Data218-1	Data219-1	Data220-1	Data221-1	Data222-1	Data223-1	GAP
x8	Master-Slave-Select-Pin-1-3	Master-Slave-Select-Pin-0-3	Selection-Ack-Pin8-1	Selection-Req-Pad1	Address-Port-1-1	Address-Port-2-1	Address-Port-3-1	Address-Port-4-1	Address-Port-5-1	Address-Port-6-1	Address-Port-7-1	Address-Port-8-1	Address-Port-9-Elite-Selected-1	RNG-Pad-0-8-1	RNG-Pad-1-8-1	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-8-1	Crossover-Out-Data-Pad-8-1	Crossover-In-Ack-Pad-8-1	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-8-1	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad8-1	SPI-Out-Line2-Pad8-1	SPI-Out-Line3-Pad8-1	SPI-Out-Line4-Pad8-1	SPI-Out-clk-Pad8-1	SPI-Out-CS-Pad8-1	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad8-4	SPI-Out-Line2-Pad8-4	SPI-Out-Line3-Pad8-4	SPI-Out-Line4-Pad8-4	SPI-Out-clk-Pad8-4	SPI-Out-CS-Pad8-4	SPI-Out-Line1-Pad8-2	SPI-Out-Line2-Pad8-2	SPI-Out-Line3-Pad8-2	SPI-Out-Line4-Pad8-2	SPI-Out-clk-Pad8-2	SPI-Out-CS-Pad8-2	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-8	PRNG-Seed-Select-Pin-1-8	PRNG-Seed-Select-Pin-2-8	PRNG-Seed-Select-Pin-3-8	Fitness-Estimation-Ack-Pin-1	Fitness-Estimation-Req1-Pad8-1	Fitness-Estimation-Req2-Pad8-1	Fitness-Estimation-Ready1-Pad8-1	Fitness-Estimation-Ready2-Pad8-1	Fitness-Estimation-Discard-Pin	Data224-1	Data225-1	Data226-1	Data227-1	Data228-1	Data229-1	Data230-1	Data231-1	Data232-1	Data233-1	Data234-1	Data235-1	Data236-1	Data237-1	Data238-1	Data239-1	Data240-1	Data241-1	Data242-1	Data243-1	Data244-1	Data245-1	Data246-1	Data247-1	Data248-1	Data249-1	Data250-1	Data251-1	Data252-1	Data253-1	Data254-1	Data255-1	GAP

x9	Master-Slave-Select-Pin-1-1	Master-Slave-Select-Pin-0-1	Selection-Req-Pad2	Selection-Ack-Pin1-2	Address-Port-1-2	Address-Port-2-2	Address-Port-3-2	Address-Port-4-2	Address-Port-5-2	Address-Port-6-2	Address-Port-7-2	Address-Port-8-2	Address-Port-9-Elite-Selected-2	RNG-Pad-0-1-2	RNG-Pad-1-1-2	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-1-2	Crossover-Out-Data-Pad-1-2	Crossover-In-Ack-Pad-1-2	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-1-2	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad1-2	SPI-Out-Line2-Pad1-2	SPI-Out-Line3-Pad1-2	SPI-Out-Line4-Pad1-2	SPI-Out-clk-Pad1-2	SPI-Out-CS-Pad1-2	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad1-1	SPI-Out-Line2-Pad1-1	SPI-Out-Line3-Pad1-1	SPI-Out-Line4-Pad1-1	SPI-Out-clk-Pad1-1	SPI-Out-CS-Pad1-1	SPI-Out-Line1-Pad1-3	SPI-Out-Line2-Pad1-3	SPI-Out-Line3-Pad1-3	SPI-Out-Line4-Pad1-3	SPI-Out-clk-Pad1-3	SPI-Out-CS-Pad1-3	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-9	PRNG-Seed-Select-Pin-1-9	PRNG-Seed-Select-Pin-2-9	PRNG-Seed-Select-Pin-3-9	Fitness-Estimation-Ack-Pin-2	Fitness-Estimation-Req1-Pad1-2	Fitness-Estimation-Req2-Pad1-2	Fitness-Estimation-Ready1-Pad1-2	Fitness-Estimation-Ready2-Pad1-2	Fitness-Estimation-Discard-Pin	Data0-2	Data1-2	Data2-2	Data3-2	Data4-2	Data5-2	Data6-2	Data7-2	Data8-2	Data9-2	Data10-2	Data11-2	Data12-2	Data13-2	Data14-2	Data15-2	Data16-2	Data17-2	Data18-2	Data19-2	Data20-2	Data21-2	Data22-2	Data23-2	Data24-2	Data25-2	Data26-2	Data27-2	Data28-2	Data29-2	Data30-2	Data31-2	GAP
x10	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin2-2	Selection-Req-Pad2	Address-Port-1-2	Address-Port-2-2	Address-Port-3-2	Address-Port-4-2	Address-Port-5-2	Address-Port-6-2	Address-Port-7-2	Address-Port-8-2	Address-Port-9-Elite-Selected-2	RNG-Pad-0-2-2	RNG-Pad-1-2-2	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-2-2	Crossover-Out-Data-Pad-2-2	Crossover-In-Ack-Pad-2-2	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-2-2	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad2-2	SPI-Out-Line2-Pad2-2	SPI-Out-Line3-Pad2-2	SPI-Out-Line4-Pad2-2	SPI-Out-clk-Pad2-2	SPI-Out-CS-Pad2-2	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad2-1	SPI-Out-Line2-Pad2-1	SPI-Out-Line3-Pad2-1	SPI-Out-Line4-Pad2-1	SPI-Out-clk-Pad2-1	SPI-Out-CS-Pad2-1	SPI-Out-Line1-Pad2-3	SPI-Out-Line2-Pad2-3	SPI-Out-Line3-Pad2-3	SPI-Out-Line4-Pad2-3	SPI-Out-clk-Pad2-3	SPI-Out-CS-Pad2-3	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-10	PRNG-Seed-Select-Pin-1-10	PRNG-Seed-Select-Pin-2-10	PRNG-Seed-Select-Pin-3-10	Fitness-Estimation-Ack-Pin-2	Fitness-Estimation-Req1-Pad2-2	Fitness-Estimation-Req2-Pad2-2	Fitness-Estimation-Ready1-Pad2-2	Fitness-Estimation-Ready2-Pad2-2	Fitness-Estimation-Discard-Pin	Data32-2	Data33-2	Data34-2	Data35-2	Data36-2	Data37-2	Data38-2	Data39-2	Data40-2	Data41-2	Data42-2	Data43-2	Data44-2	Data45-2	Data46-2	Data47-2	Data48-2	Data49-2	Data50-2	Data51-2	Data52-2	Data53-2	Data54-2	Data55-2	Data56-2	Data57-2	Data58-2	Data59-2	Data60-2	Data61-2	Data62-2	Data63-2	GAP
x11	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin3-2	Selection-Req-Pad2	Address-Port-1-2	Address-Port-2-2	Address-Port-3-2	Address-Port-4-2	Address-Port-5-2	Address-Port-6-2	Address-Port-7-2	Address-Port-8-2	Address-Port-9-Elite-Selected-2	RNG-Pad-0-3-2	RNG-Pad-1-3-2	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-3-2	Crossover-Out-Data-Pad-3-2	Crossover-In-Ack-Pad-3-2	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-3-2	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad3-2	SPI-Out-Line2-Pad3-2	SPI-Out-Line3-Pad3-2	SPI-Out-Line4-Pad3-2	SPI-Out-clk-Pad3-2	SPI-Out-CS-Pad3-2	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad3-1	SPI-Out-Line2-Pad3-1	SPI-Out-Line3-Pad3-1	SPI-Out-Line4-Pad3-1	SPI-Out-clk-Pad3-1	SPI-Out-CS-Pad3-1	SPI-Out-Line1-Pad3-3	SPI-Out-Line2-Pad3-3	SPI-Out-Line3-Pad3-3	SPI-Out-Line4-Pad3-3	SPI-Out-clk-Pad3-3	SPI-Out-CS-Pad3-3	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-11	PRNG-Seed-Select-Pin-1-11	PRNG-Seed-Select-Pin-2-11	PRNG-Seed-Select-Pin-3-11	Fitness-Estimation-Ack-Pin-2	Fitness-Estimation-Req1-Pad3-2	Fitness-Estimation-Req2-Pad3-2	Fitness-Estimation-Ready1-Pad3-2	Fitness-Estimation-Ready2-Pad3-2	Fitness-Estimation-Discard-Pin	Data64-2	Data65-2	Data66-2	Data67-2	Data68-2	Data69-2	Data70-2	Data71-2	Data72-2	Data73-2	Data74-2	Data75-2	Data76-2	Data77-2	Data78-2	Data79-2	Data80-2	Data81-2	Data82-2	Data83-2	Data84-2	Data85-2	Data86-2	Data87-2	Data88-2	Data89-2	Data90-2	Data91-2	Data92-2	Data93-2	Data94-2	Data95-2	GAP
x12	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin4-2	Selection-Req-Pad2	Address-Port-1-2	Address-Port-2-2	Address-Port-3-2	Address-Port-4-2	Address-Port-5-2	Address-Port-6-2	Address-Port-7-2	Address-Port-8-2	Address-Port-9-Elite-Selected-2	RNG-Pad-0-4-2	RNG-Pad-1-4-2	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-4-2	Crossover-Out-Data-Pad-4-2	Crossover-In-Ack-Pad-4-2	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-4-2	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad4-2	SPI-Out-Line2-Pad4-2	SPI-Out-Line3-Pad4-2	SPI-Out-Line4-Pad4-2	SPI-Out-clk-Pad4-2	SPI-Out-CS-Pad4-2	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad4-1	SPI-Out-Line2-Pad4-1	SPI-Out-Line3-Pad4-1	SPI-Out-Line4-Pad4-1	SPI-Out-clk-Pad4-1	SPI-Out-CS-Pad4-1	SPI-Out-Line1-Pad4-3	SPI-Out-Line2-Pad4-3	SPI-Out-Line3-Pad4-3	SPI-Out-Line4-Pad4-3	SPI-Out-clk-Pad4-3	SPI-Out-CS-Pad4-3	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-12	PRNG-Seed-Select-Pin-1-12	PRNG-Seed-Select-Pin-2-12	PRNG-Seed-Select-Pin-3-12	Fitness-Estimation-Ack-Pin-2	Fitness-Estimation-Req1-Pad4-2	Fitness-Estimation-Req2-Pad4-2	Fitness-Estimation-Ready1-Pad4-2	Fitness-Estimation-Ready2-Pad4-2	Fitness-Estimation-Discard-Pin	Data96-2	Data97-2	Data98-2	Data99-2	Data100-2	Data101-2	Data102-2	Data103-2	Data104-2	Data105-2	Data106-2	Data107-2	Data108-2	Data109-2	Data110-2	Data111-2	Data112-2	Data113-2	Data114-2	Data115-2	Data116-2	Data117-2	Data118-2	Data119-2	Data120-2	Data121-2	Data122-2	Data123-2	Data124-2	Data125-2	Data126-2	Data127-2	GAP
x13	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin5-2	Selection-Req-Pad2	Address-Port-1-2	Address-Port-2-2	Address-Port-3-2	Address-Port-4-2	Address-Port-5-2	Address-Port-6-2	Address-Port-7-2	Address-Port-8-2	Address-Port-9-Elite-Selected-2	RNG-Pad-0-5-2	RNG-Pad-1-5-2	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-5-2	Crossover-Out-Data-Pad-5-2	Crossover-In-Ack-Pad-5-2	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-5-2	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad5-2	SPI-Out-Line2-Pad5-2	SPI-Out-Line3-Pad5-2	SPI-Out-Line4-Pad5-2	SPI-Out-clk-Pad5-2	SPI-Out-CS-Pad5-2	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad5-1	SPI-Out-Line2-Pad5-1	SPI-Out-Line3-Pad5-1	SPI-Out-Line4-Pad5-1	SPI-Out-clk-Pad5-1	SPI-Out-CS-Pad5-1	SPI-Out-Line1-Pad5-3	SPI-Out-Line2-Pad5-3	SPI-Out-Line3-Pad5-3	SPI-Out-Line4-Pad5-3	SPI-Out-clk-Pad5-3	SPI-Out-CS-Pad5-3	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-13	PRNG-Seed-Select-Pin-1-13	PRNG-Seed-Select-Pin-2-13	PRNG-Seed-Select-Pin-3-13	Fitness-Estimation-Ack-Pin-2	Fitness-Estimation-Req1-Pad5-2	Fitness-Estimation-Req2-Pad5-2	Fitness-Estimation-Ready1-Pad5-2	Fitness-Estimation-Ready2-Pad5-2	Fitness-Estimation-Discard-Pin	Data128-2	Data129-2	Data130-2	Data131-2	Data132-2	Data133-2	Data134-2	Data135-2	Data136-2	Data137-2	Data138-2	Data139-2	Data140-2	Data141-2	Data142-2	Data143-2	Data144-2	Data145-2	Data146-2	Data147-2	Data148-2	Data149-2	Data150-2	Data151-2	Data152-2	Data153-2	Data154-2	Data155-2	Data156-2	Data157-2	Data158-2	Data159-2	GAP
x14	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin6-2	Selection-Req-Pad2	Address-Port-1-2	Address-Port-2-2	Address-Port-3-2	Address-Port-4-2	Address-Port-5-2	Address-Port-6-2	Address-Port-7-2	Address-Port-8-2	Address-Port-9-Elite-Selected-2	RNG-Pad-0-6-2	RNG-Pad-1-6-2	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-6-2	Crossover-Out-Data-Pad-6-2	Crossover-In-Ack-Pad-6-2	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-6-2	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad6-2	SPI-Out-Line2-Pad6-2	SPI-Out-Line3-Pad6-2	SPI-Out-Line4-Pad6-2	SPI-Out-clk-Pad6-2	SPI-Out-CS-Pad6-2	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad6-1	SPI-Out-Line2-Pad6-1	SPI-Out-Line3-Pad6-1	SPI-Out-Line4-Pad6-1	SPI-Out-clk-Pad6-1	SPI-Out-CS-Pad6-1	SPI-Out-Line1-Pad6-3	SPI-Out-Line2-Pad6-3	SPI-Out-Line3-Pad6-3	SPI-Out-Line4-Pad6-3	SPI-Out-clk-Pad6-3	SPI-Out-CS-Pad6-3	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-14	PRNG-Seed-Select-Pin-1-14	PRNG-Seed-Select-Pin-2-14	PRNG-Seed-Select-Pin-3-14	Fitness-Estimation-Ack-Pin-2	Fitness-Estimation-Req1-Pad6-2	Fitness-Estimation-Req2-Pad6-2	Fitness-Estimation-Ready1-Pad6-2	Fitness-Estimation-Ready2-Pad6-2	Fitness-Estimation-Discard-Pin	Data160-2	Data161-2	Data162-2	Data163-2	Data164-2	Data165-2	Data166-2	Data167-2	Data168-2	Data169-2	Data170-2	Data171-2	Data172-2	Data173-2	Data174-2	Data175-2	Data176-2	Data177-2	Data178-2	Data179-2	Data180-2	Data181-2	Data182-2	Data183-2	Data184-2	Data185-2	Data186-2	Data187-2	Data188-2	Data189-2	Data190-2	Data191-2	GAP
x15	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin7-2	Selection-Req-Pad2	Address-Port-1-2	Address-Port-2-2	Address-Port-3-2	Address-Port-4-2	Address-Port-5-2	Address-Port-6-2	Address-Port-7-2	Address-Port-8-2	Address-Port-9-Elite-Selected-2	RNG-Pad-0-7-2	RNG-Pad-1-7-2	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-7-2	Crossover-Out-Data-Pad-7-2	Crossover-In-Ack-Pad-7-2	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-7-2	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad7-2	SPI-Out-Line2-Pad7-2	SPI-Out-Line3-Pad7-2	SPI-Out-Line4-Pad7-2	SPI-Out-clk-Pad7-2	SPI-Out-CS-Pad7-2	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad7-1	SPI-Out-Line2-Pad7-1	SPI-Out-Line3-Pad7-1	SPI-Out-Line4-Pad7-1	SPI-Out-clk-Pad7-1	SPI-Out-CS-Pad7-1	SPI-Out-Line1-Pad7-3	SPI-Out-Line2-Pad7-3	SPI-Out-Line3-Pad7-3	SPI-Out-Line4-Pad7-3	SPI-Out-clk-Pad7-3	SPI-Out-CS-Pad7-3	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-15	PRNG-Seed-Select-Pin-1-15	PRNG-Seed-Select-Pin-2-15	PRNG-Seed-Select-Pin-3-15	Fitness-Estimation-Ack-Pin-2	Fitness-Estimation-Req1-Pad7-2	Fitness-Estimation-Req2-Pad7-2	Fitness-Estimation-Ready1-Pad7-2	Fitness-Estimation-Ready2-Pad7-2	Fitness-Estimation-Discard-Pin	Data192-2	Data193-2	Data194-2	Data195-2	Data196-2	Data197-2	Data198-2	Data199-2	Data200-2	Data201-2	Data202-2	Data203-2	Data204-2	Data205-2	Data206-2	Data207-2	Data208-2	Data209-2	Data210-2	Data211-2	Data212-2	Data213-2	Data214-2	Data215-2	Data216-2	Data217-2	Data218-2	Data219-2	Data220-2	Data221-2	Data222-2	Data223-2	GAP
x16	Master-Slave-Select-Pin-1-3	Master-Slave-Select-Pin-0-3	Selection-Ack-Pin8-2	Selection-Req-Pad2	Address-Port-1-2	Address-Port-2-2	Address-Port-3-2	Address-Port-4-2	Address-Port-5-2	Address-Port-6-2	Address-Port-7-2	Address-Port-8-2	Address-Port-9-Elite-Selected-2	RNG-Pad-0-8-2	RNG-Pad-1-8-2	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-8-2	Crossover-Out-Data-Pad-8-2	Crossover-In-Ack-Pad-8-2	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-8-2	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad8-2	SPI-Out-Line2-Pad8-2	SPI-Out-Line3-Pad8-2	SPI-Out-Line4-Pad8-2	SPI-Out-clk-Pad8-2	SPI-Out-CS-Pad8-2	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad8-1	SPI-Out-Line2-Pad8-1	SPI-Out-Line3-Pad8-1	SPI-Out-Line4-Pad8-1	SPI-Out-clk-Pad8-1	SPI-Out-CS-Pad8-1	SPI-Out-Line1-Pad8-3	SPI-Out-Line2-Pad8-3	SPI-Out-Line3-Pad8-3	SPI-Out-Line4-Pad8-3	SPI-Out-clk-Pad8-3	SPI-Out-CS-Pad8-3	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-16	PRNG-Seed-Select-Pin-1-16	PRNG-Seed-Select-Pin-2-16	PRNG-Seed-Select-Pin-3-16	Fitness-Estimation-Ack-Pin-2	Fitness-Estimation-Req1-Pad8-2	Fitness-Estimation-Req2-Pad8-2	Fitness-Estimation-Ready1-Pad8-2	Fitness-Estimation-Ready2-Pad8-2	Fitness-Estimation-Discard-Pin	Data224-2	Data225-2	Data226-2	Data227-2	Data228-2	Data229-2	Data230-2	Data231-2	Data232-2	Data233-2	Data234-2	Data235-2	Data236-2	Data237-2	Data238-2	Data239-2	Data240-2	Data241-2	Data242-2	Data243-2	Data244-2	Data245-2	Data246-2	Data247-2	Data248-2	Data249-2	Data250-2	Data251-2	Data252-2	Data253-2	Data254-2	Data255-2	GAP

x17	Master-Slave-Select-Pin-1-1	Master-Slave-Select-Pin-0-1	Selection-Req-Pad3	Selection-Ack-Pin1-3	Address-Port-1-3	Address-Port-2-3	Address-Port-3-3	Address-Port-4-3	Address-Port-5-3	Address-Port-6-3	Address-Port-7-3	Address-Port-8-3	Address-Port-9-Elite-Selected-3	RNG-Pad-0-1-3	RNG-Pad-1-1-3	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-1-3	Crossover-Out-Data-Pad-1-3	Crossover-In-Ack-Pad-1-3	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-1-3	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad1-3	SPI-Out-Line2-Pad1-3	SPI-Out-Line3-Pad1-3	SPI-Out-Line4-Pad1-3	SPI-Out-clk-Pad1-3	SPI-Out-CS-Pad1-3	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad1-2	SPI-Out-Line2-Pad1-2	SPI-Out-Line3-Pad1-2	SPI-Out-Line4-Pad1-2	SPI-Out-clk-Pad1-2	SPI-Out-CS-Pad1-2	SPI-Out-Line1-Pad1-4	SPI-Out-Line2-Pad1-4	SPI-Out-Line3-Pad1-4	SPI-Out-Line4-Pad1-4	SPI-Out-clk-Pad1-4	SPI-Out-CS-Pad1-4	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-8	PRNG-Seed-Select-Pin-1-8	PRNG-Seed-Select-Pin-2-8	PRNG-Seed-Select-Pin-3-8	Fitness-Estimation-Ack-Pin-3	Fitness-Estimation-Req1-Pad1-3	Fitness-Estimation-Req2-Pad1-3	Fitness-Estimation-Ready1-Pad1-3	Fitness-Estimation-Ready2-Pad1-3	Fitness-Estimation-Discard-Pin	Data0-3	Data1-3	Data2-3	Data3-3	Data4-3	Data5-3	Data6-3	Data7-3	Data8-3	Data9-3	Data10-3	Data11-3	Data12-3	Data13-3	Data14-3	Data15-3	Data16-3	Data17-3	Data18-3	Data19-3	Data20-3	Data21-3	Data22-3	Data23-3	Data24-3	Data25-3	Data26-3	Data27-3	Data28-3	Data29-3	Data30-3	Data31-3	GAP
x18	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin2-3	Selection-Req-Pad3	Address-Port-1-3	Address-Port-2-3	Address-Port-3-3	Address-Port-4-3	Address-Port-5-3	Address-Port-6-3	Address-Port-7-3	Address-Port-8-3	Address-Port-9-Elite-Selected-3	RNG-Pad-0-2-3	RNG-Pad-1-2-3	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-2-3	Crossover-Out-Data-Pad-2-3	Crossover-In-Ack-Pad-2-3	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-2-3	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad2-3	SPI-Out-Line2-Pad2-3	SPI-Out-Line3-Pad2-3	SPI-Out-Line4-Pad2-3	SPI-Out-clk-Pad2-3	SPI-Out-CS-Pad2-3	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad2-2	SPI-Out-Line2-Pad2-2	SPI-Out-Line3-Pad2-2	SPI-Out-Line4-Pad2-2	SPI-Out-clk-Pad2-2	SPI-Out-CS-Pad2-2	SPI-Out-Line1-Pad2-4	SPI-Out-Line2-Pad2-4	SPI-Out-Line3-Pad2-4	SPI-Out-Line4-Pad2-4	SPI-Out-clk-Pad2-4	SPI-Out-CS-Pad2-4	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-7	PRNG-Seed-Select-Pin-1-7	PRNG-Seed-Select-Pin-2-7	PRNG-Seed-Select-Pin-3-7	Fitness-Estimation-Ack-Pin-3	Fitness-Estimation-Req1-Pad2-3	Fitness-Estimation-Req2-Pad2-3	Fitness-Estimation-Ready1-Pad2-3	Fitness-Estimation-Ready2-Pad2-3	Fitness-Estimation-Discard-Pin	Data32-3	Data33-3	Data34-3	Data35-3	Data36-3	Data37-3	Data38-3	Data39-3	Data40-3	Data41-3	Data42-3	Data43-3	Data44-3	Data45-3	Data46-3	Data47-3	Data48-3	Data49-3	Data50-3	Data51-3	Data52-3	Data53-3	Data54-3	Data55-3	Data56-3	Data57-3	Data58-3	Data59-3	Data60-3	Data61-3	Data62-3	Data63-3	GAP
x19	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin3-3	Selection-Req-Pad3	Address-Port-1-3	Address-Port-2-3	Address-Port-3-3	Address-Port-4-3	Address-Port-5-3	Address-Port-6-3	Address-Port-7-3	Address-Port-8-3	Address-Port-9-Elite-Selected-3	RNG-Pad-0-3-3	RNG-Pad-1-3-3	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-3-3	Crossover-Out-Data-Pad-3-3	Crossover-In-Ack-Pad-3-3	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-3-3	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad3-3	SPI-Out-Line2-Pad3-3	SPI-Out-Line3-Pad3-3	SPI-Out-Line4-Pad3-3	SPI-Out-clk-Pad3-3	SPI-Out-CS-Pad3-3	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad3-2	SPI-Out-Line2-Pad3-2	SPI-Out-Line3-Pad3-2	SPI-Out-Line4-Pad3-2	SPI-Out-clk-Pad3-2	SPI-Out-CS-Pad3-2	SPI-Out-Line1-Pad3-4	SPI-Out-Line2-Pad3-4	SPI-Out-Line3-Pad3-4	SPI-Out-Line4-Pad3-4	SPI-Out-clk-Pad3-4	SPI-Out-CS-Pad3-4	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-6	PRNG-Seed-Select-Pin-1-6	PRNG-Seed-Select-Pin-2-6	PRNG-Seed-Select-Pin-3-6	Fitness-Estimation-Ack-Pin-3	Fitness-Estimation-Req1-Pad3-3	Fitness-Estimation-Req2-Pad3-3	Fitness-Estimation-Ready1-Pad3-3	Fitness-Estimation-Ready2-Pad3-3	Fitness-Estimation-Discard-Pin	Data64-3	Data65-3	Data66-3	Data67-3	Data68-3	Data69-3	Data70-3	Data71-3	Data72-3	Data73-3	Data74-3	Data75-3	Data76-3	Data77-3	Data78-3	Data79-3	Data80-3	Data81-3	Data82-3	Data83-3	Data84-3	Data85-3	Data86-3	Data87-3	Data88-3	Data89-3	Data90-3	Data91-3	Data92-3	Data93-3	Data94-3	Data95-3	GAP
x20	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin4-3	Selection-Req-Pad3	Address-Port-1-3	Address-Port-2-3	Address-Port-3-3	Address-Port-4-3	Address-Port-5-3	Address-Port-6-3	Address-Port-7-3	Address-Port-8-3	Address-Port-9-Elite-Selected-3	RNG-Pad-0-4-3	RNG-Pad-1-4-3	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-4-3	Crossover-Out-Data-Pad-4-3	Crossover-In-Ack-Pad-4-3	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-4-3	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad4-3	SPI-Out-Line2-Pad4-3	SPI-Out-Line3-Pad4-3	SPI-Out-Line4-Pad4-3	SPI-Out-clk-Pad4-3	SPI-Out-CS-Pad4-3	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad4-2	SPI-Out-Line2-Pad4-2	SPI-Out-Line3-Pad4-2	SPI-Out-Line4-Pad4-2	SPI-Out-clk-Pad4-2	SPI-Out-CS-Pad4-2	SPI-Out-Line1-Pad4-4	SPI-Out-Line2-Pad4-4	SPI-Out-Line3-Pad4-4	SPI-Out-Line4-Pad4-4	SPI-Out-clk-Pad4-4	SPI-Out-CS-Pad4-4	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-5	PRNG-Seed-Select-Pin-1-5	PRNG-Seed-Select-Pin-2-5	PRNG-Seed-Select-Pin-3-5	Fitness-Estimation-Ack-Pin-3	Fitness-Estimation-Req1-Pad4-3	Fitness-Estimation-Req2-Pad4-3	Fitness-Estimation-Ready1-Pad4-3	Fitness-Estimation-Ready2-Pad4-3	Fitness-Estimation-Discard-Pin	Data96-3	Data97-3	Data98-3	Data99-3	Data100-3	Data101-3	Data102-3	Data103-3	Data104-3	Data105-3	Data106-3	Data107-3	Data108-3	Data109-3	Data110-3	Data111-3	Data112-3	Data113-3	Data114-3	Data115-3	Data116-3	Data117-3	Data118-3	Data119-3	Data120-3	Data121-3	Data122-3	Data123-3	Data124-3	Data125-3	Data126-3	Data127-3	GAP
x21	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin5-3	Selection-Req-Pad3	Address-Port-1-3	Address-Port-2-3	Address-Port-3-3	Address-Port-4-3	Address-Port-5-3	Address-Port-6-3	Address-Port-7-3	Address-Port-8-3	Address-Port-9-Elite-Selected-3	RNG-Pad-0-5-3	RNG-Pad-1-5-3	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-5-3	Crossover-Out-Data-Pad-5-3	Crossover-In-Ack-Pad-5-3	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-5-3	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad5-3	SPI-Out-Line2-Pad5-3	SPI-Out-Line3-Pad5-3	SPI-Out-Line4-Pad5-3	SPI-Out-clk-Pad5-3	SPI-Out-CS-Pad5-3	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad5-2	SPI-Out-Line2-Pad5-2	SPI-Out-Line3-Pad5-2	SPI-Out-Line4-Pad5-2	SPI-Out-clk-Pad5-2	SPI-Out-CS-Pad5-2	SPI-Out-Line1-Pad5-4	SPI-Out-Line2-Pad5-4	SPI-Out-Line3-Pad5-4	SPI-Out-Line4-Pad5-4	SPI-Out-clk-Pad5-4	SPI-Out-CS-Pad5-4	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-4	PRNG-Seed-Select-Pin-1-4	PRNG-Seed-Select-Pin-2-4	PRNG-Seed-Select-Pin-3-4	Fitness-Estimation-Ack-Pin-3	Fitness-Estimation-Req1-Pad5-3	Fitness-Estimation-Req2-Pad5-3	Fitness-Estimation-Ready1-Pad5-3	Fitness-Estimation-Ready2-Pad5-3	Fitness-Estimation-Discard-Pin	Data128-3	Data129-3	Data130-3	Data131-3	Data132-3	Data133-3	Data134-3	Data135-3	Data136-3	Data137-3	Data138-3	Data139-3	Data140-3	Data141-3	Data142-3	Data143-3	Data144-3	Data145-3	Data146-3	Data147-3	Data148-3	Data149-3	Data150-3	Data151-3	Data152-3	Data153-3	Data154-3	Data155-3	Data156-3	Data157-3	Data158-3	Data159-3	GAP
x22	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin6-3	Selection-Req-Pad3	Address-Port-1-3	Address-Port-2-3	Address-Port-3-3	Address-Port-4-3	Address-Port-5-3	Address-Port-6-3	Address-Port-7-3	Address-Port-8-3	Address-Port-9-Elite-Selected-3	RNG-Pad-0-6-3	RNG-Pad-1-6-3	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-6-3	Crossover-Out-Data-Pad-6-3	Crossover-In-Ack-Pad-6-3	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-6-3	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad6-3	SPI-Out-Line2-Pad6-3	SPI-Out-Line3-Pad6-3	SPI-Out-Line4-Pad6-3	SPI-Out-clk-Pad6-3	SPI-Out-CS-Pad6-3	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad6-2	SPI-Out-Line2-Pad6-2	SPI-Out-Line3-Pad6-2	SPI-Out-Line4-Pad6-2	SPI-Out-clk-Pad6-2	SPI-Out-CS-Pad6-2	SPI-Out-Line1-Pad6-4	SPI-Out-Line2-Pad6-4	SPI-Out-Line3-Pad6-4	SPI-Out-Line4-Pad6-4	SPI-Out-clk-Pad6-4	SPI-Out-CS-Pad6-4	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-3	PRNG-Seed-Select-Pin-1-3	PRNG-Seed-Select-Pin-2-3	PRNG-Seed-Select-Pin-3-3	Fitness-Estimation-Ack-Pin-3	Fitness-Estimation-Req1-Pad6-3	Fitness-Estimation-Req2-Pad6-3	Fitness-Estimation-Ready1-Pad6-3	Fitness-Estimation-Ready2-Pad6-3	Fitness-Estimation-Discard-Pin	Data160-3	Data161-3	Data162-3	Data163-3	Data164-3	Data165-3	Data166-3	Data167-3	Data168-3	Data169-3	Data170-3	Data171-3	Data172-3	Data173-3	Data174-3	Data175-3	Data176-3	Data177-3	Data178-3	Data179-3	Data180-3	Data181-3	Data182-3	Data183-3	Data184-3	Data185-3	Data186-3	Data187-3	Data188-3	Data189-3	Data190-3	Data191-3	GAP
x23	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin7-3	Selection-Req-Pad3	Address-Port-1-3	Address-Port-2-3	Address-Port-3-3	Address-Port-4-3	Address-Port-5-3	Address-Port-6-3	Address-Port-7-3	Address-Port-8-3	Address-Port-9-Elite-Selected-3	RNG-Pad-0-7-3	RNG-Pad-1-7-3	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-7-3	Crossover-Out-Data-Pad-7-3	Crossover-In-Ack-Pad-7-3	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-7-3	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad7-3	SPI-Out-Line2-Pad7-3	SPI-Out-Line3-Pad7-3	SPI-Out-Line4-Pad7-3	SPI-Out-clk-Pad7-3	SPI-Out-CS-Pad7-3	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad7-2	SPI-Out-Line2-Pad7-2	SPI-Out-Line3-Pad7-2	SPI-Out-Line4-Pad7-2	SPI-Out-clk-Pad7-2	SPI-Out-CS-Pad7-2	SPI-Out-Line1-Pad7-4	SPI-Out-Line2-Pad7-4	SPI-Out-Line3-Pad7-4	SPI-Out-Line4-Pad7-4	SPI-Out-clk-Pad7-4	SPI-Out-CS-Pad7-4	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-2	PRNG-Seed-Select-Pin-1-2	PRNG-Seed-Select-Pin-2-2	PRNG-Seed-Select-Pin-3-2	Fitness-Estimation-Ack-Pin-3	Fitness-Estimation-Req1-Pad7-3	Fitness-Estimation-Req2-Pad7-3	Fitness-Estimation-Ready1-Pad7-3	Fitness-Estimation-Ready2-Pad7-3	Fitness-Estimation-Discard-Pin	Data192-3	Data193-3	Data194-3	Data195-3	Data196-3	Data197-3	Data198-3	Data199-3	Data200-3	Data201-3	Data202-3	Data203-3	Data204-3	Data205-3	Data206-3	Data207-3	Data208-3	Data209-3	Data210-3	Data211-3	Data212-3	Data213-3	Data214-3	Data215-3	Data216-3	Data217-3	Data218-3	Data219-3	Data220-3	Data221-3	Data222-3	Data223-3	GAP
x24	Master-Slave-Select-Pin-1-3	Master-Slave-Select-Pin-0-3	Selection-Ack-Pin8-3	Selection-Req-Pad3	Address-Port-1-3	Address-Port-2-3	Address-Port-3-3	Address-Port-4-3	Address-Port-5-3	Address-Port-6-3	Address-Port-7-3	Address-Port-8-3	Address-Port-9-Elite-Selected-3	RNG-Pad-0-8-3	RNG-Pad-1-8-3	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-8-3	Crossover-Out-Data-Pad-8-3	Crossover-In-Ack-Pad-8-3	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-8-3	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad8-3	SPI-Out-Line2-Pad8-3	SPI-Out-Line3-Pad8-3	SPI-Out-Line4-Pad8-3	SPI-Out-clk-Pad8-3	SPI-Out-CS-Pad8-3	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad8-2	SPI-Out-Line2-Pad8-2	SPI-Out-Line3-Pad8-2	SPI-Out-Line4-Pad8-2	SPI-Out-clk-Pad8-2	SPI-Out-CS-Pad8-2	SPI-Out-Line1-Pad8-4	SPI-Out-Line2-Pad8-4	SPI-Out-Line3-Pad8-4	SPI-Out-Line4-Pad8-4	SPI-Out-clk-Pad8-4	SPI-Out-CS-Pad8-4	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-1	PRNG-Seed-Select-Pin-1-1	PRNG-Seed-Select-Pin-2-1	PRNG-Seed-Select-Pin-3-1	Fitness-Estimation-Ack-Pin-3	Fitness-Estimation-Req1-Pad8-3	Fitness-Estimation-Req2-Pad8-3	Fitness-Estimation-Ready1-Pad8-3	Fitness-Estimation-Ready2-Pad8-3	Fitness-Estimation-Discard-Pin	Data224-3	Data225-3	Data226-3	Data227-3	Data228-3	Data229-3	Data230-3	Data231-3	Data232-3	Data233-3	Data234-3	Data235-3	Data236-3	Data237-3	Data238-3	Data239-3	Data240-3	Data241-3	Data242-3	Data243-3	Data244-3	Data245-3	Data246-3	Data247-3	Data248-3	Data249-3	Data250-3	Data251-3	Data252-3	Data253-3	Data254-3	Data255-3	GAP

x25	Master-Slave-Select-Pin-1-1	Master-Slave-Select-Pin-0-1	Selection-Req-Pad4	Selection-Ack-Pin1-4	Address-Port-1-4	Address-Port-2-4	Address-Port-3-4	Address-Port-4-4	Address-Port-5-4	Address-Port-6-4	Address-Port-7-4	Address-Port-8-4	Address-Port-9-Elite-Selected-4	RNG-Pad-0-1-4	RNG-Pad-1-1-4	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-1-4	Crossover-Out-Data-Pad-1-4	Crossover-In-Ack-Pad-1-4	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-1-4	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad1-4	SPI-Out-Line2-Pad1-4	SPI-Out-Line3-Pad1-4	SPI-Out-Line4-Pad1-4	SPI-Out-clk-Pad1-4	SPI-Out-CS-Pad1-4	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad1-3	SPI-Out-Line2-Pad1-3	SPI-Out-Line3-Pad1-3	SPI-Out-Line4-Pad1-3	SPI-Out-clk-Pad1-3	SPI-Out-CS-Pad1-3	SPI-Out-Line1-Pad1-1	SPI-Out-Line2-Pad1-1	SPI-Out-Line3-Pad1-1	SPI-Out-Line4-Pad1-1	SPI-Out-clk-Pad1-1	SPI-Out-CS-Pad1-1	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-16	PRNG-Seed-Select-Pin-1-16	PRNG-Seed-Select-Pin-2-16	PRNG-Seed-Select-Pin-3-16	Fitness-Estimation-Ack-Pin-4	Fitness-Estimation-Req1-Pad1-4	Fitness-Estimation-Req2-Pad1-4	Fitness-Estimation-Ready1-Pad1-4	Fitness-Estimation-Ready2-Pad1-4	Fitness-Estimation-Discard-Pin	Data0-4	Data1-4	Data2-4	Data3-4	Data4-4	Data5-4	Data6-4	Data7-4	Data8-4	Data9-4	Data10-4	Data11-4	Data12-4	Data13-4	Data14-4	Data15-4	Data16-4	Data17-4	Data18-4	Data19-4	Data20-4	Data21-4	Data22-4	Data23-4	Data24-4	Data25-4	Data26-4	Data27-4	Data28-4	Data29-4	Data30-4	Data31-4	GAP
x26	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin2-4	Selection-Req-Pad4	Address-Port-1-4	Address-Port-2-4	Address-Port-3-4	Address-Port-4-4	Address-Port-5-4	Address-Port-6-4	Address-Port-7-4	Address-Port-8-4	Address-Port-9-Elite-Selected-4	RNG-Pad-0-2-4	RNG-Pad-1-2-4	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-2-4	Crossover-Out-Data-Pad-2-4	Crossover-In-Ack-Pad-2-4	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-2-4	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad2-4	SPI-Out-Line2-Pad2-4	SPI-Out-Line3-Pad2-4	SPI-Out-Line4-Pad2-4	SPI-Out-clk-Pad2-4	SPI-Out-CS-Pad2-4	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad2-3	SPI-Out-Line2-Pad2-3	SPI-Out-Line3-Pad2-3	SPI-Out-Line4-Pad2-3	SPI-Out-clk-Pad2-3	SPI-Out-CS-Pad2-3	SPI-Out-Line1-Pad2-1	SPI-Out-Line2-Pad2-1	SPI-Out-Line3-Pad2-1	SPI-Out-Line4-Pad2-1	SPI-Out-clk-Pad2-1	SPI-Out-CS-Pad2-1	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-15	PRNG-Seed-Select-Pin-1-15	PRNG-Seed-Select-Pin-2-15	PRNG-Seed-Select-Pin-3-15	Fitness-Estimation-Ack-Pin-4	Fitness-Estimation-Req1-Pad2-4	Fitness-Estimation-Req2-Pad2-4	Fitness-Estimation-Ready1-Pad2-4	Fitness-Estimation-Ready2-Pad2-4	Fitness-Estimation-Discard-Pin	Data32-4	Data33-4	Data34-4	Data35-4	Data36-4	Data37-4	Data38-4	Data39-4	Data40-4	Data41-4	Data42-4	Data43-4	Data44-4	Data45-4	Data46-4	Data47-4	Data48-4	Data49-4	Data50-4	Data51-4	Data52-4	Data53-4	Data54-4	Data55-4	Data56-4	Data57-4	Data58-4	Data59-4	Data60-4	Data61-4	Data62-4	Data63-4	GAP
x27	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin3-4	Selection-Req-Pad4	Address-Port-1-4	Address-Port-2-4	Address-Port-3-4	Address-Port-4-4	Address-Port-5-4	Address-Port-6-4	Address-Port-7-4	Address-Port-8-4	Address-Port-9-Elite-Selected-4	RNG-Pad-0-3-4	RNG-Pad-1-3-4	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-3-4	Crossover-Out-Data-Pad-3-4	Crossover-In-Ack-Pad-3-4	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-3-4	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad3-4	SPI-Out-Line2-Pad3-4	SPI-Out-Line3-Pad3-4	SPI-Out-Line4-Pad3-4	SPI-Out-clk-Pad3-4	SPI-Out-CS-Pad3-4	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad3-3	SPI-Out-Line2-Pad3-3	SPI-Out-Line3-Pad3-3	SPI-Out-Line4-Pad3-3	SPI-Out-clk-Pad3-3	SPI-Out-CS-Pad3-3	SPI-Out-Line1-Pad3-1	SPI-Out-Line2-Pad3-1	SPI-Out-Line3-Pad3-1	SPI-Out-Line4-Pad3-1	SPI-Out-clk-Pad3-1	SPI-Out-CS-Pad3-1	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-14	PRNG-Seed-Select-Pin-1-14	PRNG-Seed-Select-Pin-2-14	PRNG-Seed-Select-Pin-3-14	Fitness-Estimation-Ack-Pin-4	Fitness-Estimation-Req1-Pad3-4	Fitness-Estimation-Req2-Pad3-4	Fitness-Estimation-Ready1-Pad3-4	Fitness-Estimation-Ready2-Pad3-4	Fitness-Estimation-Discard-Pin	Data64-4	Data65-4	Data66-4	Data67-4	Data68-4	Data69-4	Data70-4	Data71-4	Data72-4	Data73-4	Data74-4	Data75-4	Data76-4	Data77-4	Data78-4	Data79-4	Data80-4	Data81-4	Data82-4	Data83-4	Data84-4	Data85-4	Data86-4	Data87-4	Data88-4	Data89-4	Data90-4	Data91-4	Data92-4	Data93-4	Data94-4	Data95-4	GAP
x28	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin4-4	Selection-Req-Pad4	Address-Port-1-4	Address-Port-2-4	Address-Port-3-4	Address-Port-4-4	Address-Port-5-4	Address-Port-6-4	Address-Port-7-4	Address-Port-8-4	Address-Port-9-Elite-Selected-4	RNG-Pad-0-4-4	RNG-Pad-1-4-4	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-4-4	Crossover-Out-Data-Pad-4-4	Crossover-In-Ack-Pad-4-4	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-4-4	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad4-4	SPI-Out-Line2-Pad4-4	SPI-Out-Line3-Pad4-4	SPI-Out-Line4-Pad4-4	SPI-Out-clk-Pad4-4	SPI-Out-CS-Pad4-4	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad4-3	SPI-Out-Line2-Pad4-3	SPI-Out-Line3-Pad4-3	SPI-Out-Line4-Pad4-3	SPI-Out-clk-Pad4-3	SPI-Out-CS-Pad4-3	SPI-Out-Line1-Pad4-1	SPI-Out-Line2-Pad4-1	SPI-Out-Line3-Pad4-1	SPI-Out-Line4-Pad4-1	SPI-Out-clk-Pad4-1	SPI-Out-CS-Pad4-1	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-13	PRNG-Seed-Select-Pin-1-13	PRNG-Seed-Select-Pin-2-13	PRNG-Seed-Select-Pin-3-13	Fitness-Estimation-Ack-Pin-4	Fitness-Estimation-Req1-Pad4-4	Fitness-Estimation-Req2-Pad4-4	Fitness-Estimation-Ready1-Pad4-4	Fitness-Estimation-Ready2-Pad4-4	Fitness-Estimation-Discard-Pin	Data96-4	Data97-4	Data98-4	Data99-4	Data100-4	Data101-4	Data102-4	Data103-4	Data104-4	Data105-4	Data106-4	Data107-4	Data108-4	Data109-4	Data110-4	Data111-4	Data112-4	Data113-4	Data114-4	Data115-4	Data116-4	Data117-4	Data118-4	Data119-4	Data120-4	Data121-4	Data122-4	Data123-4	Data124-4	Data125-4	Data126-4	Data127-4	GAP
x29	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin5-4	Selection-Req-Pad4	Address-Port-1-4	Address-Port-2-4	Address-Port-3-4	Address-Port-4-4	Address-Port-5-4	Address-Port-6-4	Address-Port-7-4	Address-Port-8-4	Address-Port-9-Elite-Selected-4	RNG-Pad-0-5-4	RNG-Pad-1-5-4	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-5-4	Crossover-Out-Data-Pad-5-4	Crossover-In-Ack-Pad-5-4	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-5-4	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad5-4	SPI-Out-Line2-Pad5-4	SPI-Out-Line3-Pad5-4	SPI-Out-Line4-Pad5-4	SPI-Out-clk-Pad5-4	SPI-Out-CS-Pad5-4	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad5-3	SPI-Out-Line2-Pad5-3	SPI-Out-Line3-Pad5-3	SPI-Out-Line4-Pad5-3	SPI-Out-clk-Pad5-3	SPI-Out-CS-Pad5-3	SPI-Out-Line1-Pad5-1	SPI-Out-Line2-Pad5-1	SPI-Out-Line3-Pad5-1	SPI-Out-Line4-Pad5-1	SPI-Out-clk-Pad5-1	SPI-Out-CS-Pad5-1	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-12	PRNG-Seed-Select-Pin-1-12	PRNG-Seed-Select-Pin-2-12	PRNG-Seed-Select-Pin-3-12	Fitness-Estimation-Ack-Pin-4	Fitness-Estimation-Req1-Pad5-4	Fitness-Estimation-Req2-Pad5-4	Fitness-Estimation-Ready1-Pad5-4	Fitness-Estimation-Ready2-Pad5-4	Fitness-Estimation-Discard-Pin	Data128-4	Data129-4	Data130-4	Data131-4	Data132-4	Data133-4	Data134-4	Data135-4	Data136-4	Data137-4	Data138-4	Data139-4	Data140-4	Data141-4	Data142-4	Data143-4	Data144-4	Data145-4	Data146-4	Data147-4	Data148-4	Data149-4	Data150-4	Data151-4	Data152-4	Data153-4	Data154-4	Data155-4	Data156-4	Data157-4	Data158-4	Data159-4	GAP
x30	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin6-4	Selection-Req-Pad4	Address-Port-1-4	Address-Port-2-4	Address-Port-3-4	Address-Port-4-4	Address-Port-5-4	Address-Port-6-4	Address-Port-7-4	Address-Port-8-4	Address-Port-9-Elite-Selected-4	RNG-Pad-0-6-4	RNG-Pad-1-6-4	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-6-4	Crossover-Out-Data-Pad-6-4	Crossover-In-Ack-Pad-6-4	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-6-4	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad6-4	SPI-Out-Line2-Pad6-4	SPI-Out-Line3-Pad6-4	SPI-Out-Line4-Pad6-4	SPI-Out-clk-Pad6-4	SPI-Out-CS-Pad6-4	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad6-3	SPI-Out-Line2-Pad6-3	SPI-Out-Line3-Pad6-3	SPI-Out-Line4-Pad6-3	SPI-Out-clk-Pad6-3	SPI-Out-CS-Pad6-3	SPI-Out-Line1-Pad6-1	SPI-Out-Line2-Pad6-1	SPI-Out-Line3-Pad6-1	SPI-Out-Line4-Pad6-1	SPI-Out-clk-Pad6-1	SPI-Out-CS-Pad6-1	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-11	PRNG-Seed-Select-Pin-1-11	PRNG-Seed-Select-Pin-2-11	PRNG-Seed-Select-Pin-3-11	Fitness-Estimation-Ack-Pin-4	Fitness-Estimation-Req1-Pad6-4	Fitness-Estimation-Req2-Pad6-4	Fitness-Estimation-Ready1-Pad6-4	Fitness-Estimation-Ready2-Pad6-4	Fitness-Estimation-Discard-Pin	Data160-4	Data161-4	Data162-4	Data163-4	Data164-4	Data165-4	Data166-4	Data167-4	Data168-4	Data169-4	Data170-4	Data171-4	Data172-4	Data173-4	Data174-4	Data175-4	Data176-4	Data177-4	Data178-4	Data179-4	Data180-4	Data181-4	Data182-4	Data183-4	Data184-4	Data185-4	Data186-4	Data187-4	Data188-4	Data189-4	Data190-4	Data191-4	GAP
x31	Master-Slave-Select-Pin-1-2	Master-Slave-Select-Pin-0-2	Selection-Ack-Pin7-4	Selection-Req-Pad4	Address-Port-1-4	Address-Port-2-4	Address-Port-3-4	Address-Port-4-4	Address-Port-5-4	Address-Port-6-4	Address-Port-7-4	Address-Port-8-4	Address-Port-9-Elite-Selected-4	RNG-Pad-0-7-4	RNG-Pad-1-7-4	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-7-4	Crossover-Out-Data-Pad-7-4	Crossover-In-Ack-Pad-7-4	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-7-4	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad7-4	SPI-Out-Line2-Pad7-4	SPI-Out-Line3-Pad7-4	SPI-Out-Line4-Pad7-4	SPI-Out-clk-Pad7-4	SPI-Out-CS-Pad7-4	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad7-3	SPI-Out-Line2-Pad7-3	SPI-Out-Line3-Pad7-3	SPI-Out-Line4-Pad7-3	SPI-Out-clk-Pad7-3	SPI-Out-CS-Pad7-3	SPI-Out-Line1-Pad7-1	SPI-Out-Line2-Pad7-1	SPI-Out-Line3-Pad7-1	SPI-Out-Line4-Pad7-1	SPI-Out-clk-Pad7-1	SPI-Out-CS-Pad7-1	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-10	PRNG-Seed-Select-Pin-1-10	PRNG-Seed-Select-Pin-2-10	PRNG-Seed-Select-Pin-3-10	Fitness-Estimation-Ack-Pin-4	Fitness-Estimation-Req1-Pad7-4	Fitness-Estimation-Req2-Pad7-4	Fitness-Estimation-Ready1-Pad7-4	Fitness-Estimation-Ready2-Pad7-4	Fitness-Estimation-Discard-Pin	Data192-4	Data193-4	Data194-4	Data195-4	Data196-4	Data197-4	Data198-4	Data199-4	Data200-4	Data201-4	Data202-4	Data203-4	Data204-4	Data205-4	Data206-4	Data207-4	Data208-4	Data209-4	Data210-4	Data211-4	Data212-4	Data213-4	Data214-4	Data215-4	Data216-4	Data217-4	Data218-4	Data219-4	Data220-4	Data221-4	Data222-4	Data223-4	GAP
x32	Master-Slave-Select-Pin-1-3	Master-Slave-Select-Pin-0-3	Selection-Ack-Pin8-4	Selection-Req-Pad4	Address-Port-1-4	Address-Port-2-4	Address-Port-3-4	Address-Port-4-4	Address-Port-5-4	Address-Port-6-4	Address-Port-7-4	Address-Port-8-4	Address-Port-9-Elite-Selected-4	RNG-Pad-0-8-4	RNG-Pad-1-8-4	Crossover-Out-Ack-Pin	Crossover-Out-Req-Pad-8-4	Crossover-Out-Data-Pad-8-4	Crossover-In-Ack-Pad-8-4	Crossover-In-Req-Pin	Crossover-In-Data-Pin	Chromosome-Resolution-Pin	Fitness-Resolution-Pin	Best-Found-Emmigration-Pin	No-Elitism-Pin	Dual-Ram-Pin	Data-Ready-Pad-8-4	Restart-Pin	Stop-Pin	Clock-1-Pin	Clock-2-Pin	Population-Size-Pin-0	Population-Size-Pin-1	Random-Immigrants-Gap-Pin-1	Random-Immigrants-Gap-Pin-0	Mutation-Rate-Pin-0	Mutation-Rate-Pin-1	Mutation-Rate-Pin-2	Mutation-Rate-Pin-3	Mutation-Rate-Pin-4	Mutation-Rate-Pin-5	Mutation-Rate-Pin-6	Crossover-Rate-Pin-0	Crossover-Rate-Pin-1	Crossover-Rate-Pin-2	Crossover-Rate-Pin-3	Crossover-Rate-Pin-4	Crossover-Rate-Pin-5	Crossover-Rate-Pin-6	Migration-Gap-Pin-1	Migration-Gap-Pin-0	SPI-Out-Line1-Pad8-4	SPI-Out-Line2-Pad8-4	SPI-Out-Line3-Pad8-4	SPI-Out-Line4-Pad8-4	SPI-Out-clk-Pad8-4	SPI-Out-CS-Pad8-4	Second-SPI-Ready-Pin	SPI-Out-Line1-Pad8-3	SPI-Out-Line2-Pad8-3	SPI-Out-Line3-Pad8-3	SPI-Out-Line4-Pad8-3	SPI-Out-clk-Pad8-3	SPI-Out-CS-Pad8-3	SPI-Out-Line1-Pad8-1	SPI-Out-Line2-Pad8-1	SPI-Out-Line3-Pad8-1	SPI-Out-Line4-Pad8-1	SPI-Out-clk-Pad8-1	SPI-Out-CS-Pad8-1	Fitness-or-Cost-Pin	Tournament-Size-Pin-1	Tournament-Size-Pin-0	Iteration-Number-Pin-0	Iteration-Number-Pin-1	Iteration-Number-Pin-2	Uniform-Mutation-Pin	One-Point-Mutation-Pin	Uniform-Crossover-Pin	Crossover-Type-Pin-1	Crossover-Type-Pin-0	Pipeline-Stages-Pin-3	Pipeline-Stages-Pin-2	Pipeline-Stages-Pin-1	Pipeline-Stages-Pin-0	PRNG-Seed-Select-Pin-0-9	PRNG-Seed-Select-Pin-1-9	PRNG-Seed-Select-Pin-2-9	PRNG-Seed-Select-Pin-3-9	Fitness-Estimation-Ack-Pin-4	Fitness-Estimation-Req1-Pad8-4	Fitness-Estimation-Req2-Pad8-4	Fitness-Estimation-Ready1-Pad8-4	Fitness-Estimation-Ready2-Pad8-4	Fitness-Estimation-Discard-Pin	Data224-4	Data225-4	Data226-4	Data227-4	Data228-4	Data229-4	Data230-4	Data231-4	Data232-4	Data233-4	Data234-4	Data235-4	Data236-4	Data237-4	Data238-4	Data239-4	Data240-4	Data241-4	Data242-4	Data243-4	Data244-4	Data245-4	Data246-4	Data247-4	Data248-4	Data249-4	Data250-4	Data251-4	Data252-4	Data253-4	Data254-4	Data255-4	GAP
	

*Fitness Computation Units
x33	Req1-1	Ready1-1	Fitness-Estimation-Ack-Pin1-1 DData0-1 DData1-1 DData2-1 DData3-1 DData4-1 DData5-1 DData6-1 DData7-1 DData8-1 DData9-1 DData10-1 DData11-1 DData12-1 DData13-1 DData14-1 DData15-1 Data16-1 Data17-1 Data18-1 Data19-1 Data20-1 Data21-1 Data22-1 Data23-1 Data24-1 Data25-1 Data26-1 Data27-1 Data28-1 Data29-1 Data30-1 Data31-1 DData32-1 DData33-1 DData34-1 DData35-1 DData36-1 DData37-1 DData38-1 DData39-1 DData40-1 DData41-1 DData42-1 DData43-1 DData44-1 DData45-1 DData46-1 DData47-1 Data48-1 Data49-1 Data50-1 Data51-1 Data52-1 Data53-1 Data54-1 Data55-1 Data56-1 Data57-1 Data58-1 Data59-1 Data60-1 Data61-1 Data62-1 Data63-1 DData64-1 DData65-1 DData66-1 DData67-1 DData68-1 DData69-1 DData70-1 DData71-1 DData72-1 DData73-1 DData74-1 DData75-1 DData76-1 DData77-1 DData78-1 DData79-1 Data80-1 Data81-1 Data82-1 Data83-1 Data84-1 Data85-1 Data86-1 Data87-1 Data88-1 Data89-1 Data90-1 Data91-1 Data92-1 Data93-1 Data94-1 Data95-1 DData96-1 DData97-1 DData98-1 DData99-1 DData100-1 DData101-1 DData102-1 DData103-1 DData104-1 DData105-1 DData106-1 DData107-1 DData108-1 DData109-1 DData110-1 DData111-1 Data112-1 Data113-1 Data114-1 Data115-1 Data116-1 Data117-1 Data118-1 Data119-1 Data120-1 Data121-1 Data122-1 Data123-1 Data124-1 Data125-1 Data126-1 Data127-1 DData128-1 DData129-1 DData130-1 DData131-1 DData132-1 DData133-1 DData134-1 DData135-1 DData136-1 DData137-1 DData138-1 DData139-1 DData140-1 DData141-1 DData142-1 DData143-1 Data144-1 Data145-1 Data146-1 Data147-1 Data148-1 Data149-1 Data150-1 Data151-1 Data152-1 Data153-1 Data154-1 Data155-1 Data156-1 Data157-1 Data158-1 Data159-1 DData160-1 DData161-1 DData162-1 DData163-1 DData164-1 DData165-1 DData166-1 DData167-1 DData168-1 DData169-1 DData170-1 DData171-1 DData172-1 DData173-1 DData174-1 DData175-1 Data176-1 Data177-1 Data178-1 Data179-1 Data180-1 Data181-1 Data182-1 Data183-1 Data184-1 Data185-1 Data186-1 Data187-1 Data188-1 Data189-1 Data190-1 Data191-1 DData192-1 DData193-1 DData194-1 DData195-1 DData196-1 DData197-1 DData198-1 DData199-1 DData200-1 DData201-1 DData202-1 DData203-1 DData204-1 DData205-1 DData206-1 DData207-1 Data208-1 Data209-1 Data210-1 Data211-1 Data212-1 Data213-1 Data214-1 Data215-1 Data216-1 Data217-1 Data218-1 Data219-1 Data220-1 Data221-1 Data222-1 Data223-1 DData224-1 DData225-1 DData226-1 DData227-1 DData228-1 DData229-1 DData230-1 DData231-1 DData232-1 DData233-1 DData234-1 DData235-1 DData236-1 DData237-1 DData238-1 DData239-1 Data240-1 Data241-1 Data242-1 Data243-1 Data244-1 Data245-1 Data246-1 Data247-1 Data248-1 Data249-1 Data250-1 Data251-1 Data252-1 Data253-1 Data254-1 Data255-1 Out0-1-1 Out1-1-1 Out2-1-1 Out3-1-1 Out4-1-1 Out5-1-1 Out6-1-1 Out7-1-1 Out8-1-1	RoyalRoad
x34	Req2-1	Ready2-1	Fitness-Estimation-Ack-Pin2-1 DData0-1 DData1-1 DData2-1 DData3-1 DData4-1 DData5-1 DData6-1 DData7-1 DData8-1 DData9-1 DData10-1 DData11-1 DData12-1 DData13-1 DData14-1 DData15-1 Data16-1 Data17-1 Data18-1 Data19-1 Data20-1 Data21-1 Data22-1 Data23-1 Data24-1 Data25-1 Data26-1 Data27-1 Data28-1 Data29-1 Data30-1 Data31-1 DData32-1 DData33-1 DData34-1 DData35-1 DData36-1 DData37-1 DData38-1 DData39-1 DData40-1 DData41-1 DData42-1 DData43-1 DData44-1 DData45-1 DData46-1 DData47-1 Data48-1 Data49-1 Data50-1 Data51-1 Data52-1 Data53-1 Data54-1 Data55-1 Data56-1 Data57-1 Data58-1 Data59-1 Data60-1 Data61-1 Data62-1 Data63-1 DData64-1 DData65-1 DData66-1 DData67-1 DData68-1 DData69-1 DData70-1 DData71-1 DData72-1 DData73-1 DData74-1 DData75-1 DData76-1 DData77-1 DData78-1 DData79-1 Data80-1 Data81-1 Data82-1 Data83-1 Data84-1 Data85-1 Data86-1 Data87-1 Data88-1 Data89-1 Data90-1 Data91-1 Data92-1 Data93-1 Data94-1 Data95-1 DData96-1 DData97-1 DData98-1 DData99-1 DData100-1 DData101-1 DData102-1 DData103-1 DData104-1 DData105-1 DData106-1 DData107-1 DData108-1 DData109-1 DData110-1 DData111-1 Data112-1 Data113-1 Data114-1 Data115-1 Data116-1 Data117-1 Data118-1 Data119-1 Data120-1 Data121-1 Data122-1 Data123-1 Data124-1 Data125-1 Data126-1 Data127-1 DData128-1 DData129-1 DData130-1 DData131-1 DData132-1 DData133-1 DData134-1 DData135-1 DData136-1 DData137-1 DData138-1 DData139-1 DData140-1 DData141-1 DData142-1 DData143-1 Data144-1 Data145-1 Data146-1 Data147-1 Data148-1 Data149-1 Data150-1 Data151-1 Data152-1 Data153-1 Data154-1 Data155-1 Data156-1 Data157-1 Data158-1 Data159-1 DData160-1 DData161-1 DData162-1 DData163-1 DData164-1 DData165-1 DData166-1 DData167-1 DData168-1 DData169-1 DData170-1 DData171-1 DData172-1 DData173-1 DData174-1 DData175-1 Data176-1 Data177-1 Data178-1 Data179-1 Data180-1 Data181-1 Data182-1 Data183-1 Data184-1 Data185-1 Data186-1 Data187-1 Data188-1 Data189-1 Data190-1 Data191-1 DData192-1 DData193-1 DData194-1 DData195-1 DData196-1 DData197-1 DData198-1 DData199-1 DData200-1 DData201-1 DData202-1 DData203-1 DData204-1 DData205-1 DData206-1 DData207-1 Data208-1 Data209-1 Data210-1 Data211-1 Data212-1 Data213-1 Data214-1 Data215-1 Data216-1 Data217-1 Data218-1 Data219-1 Data220-1 Data221-1 Data222-1 Data223-1 DData224-1 DData225-1 DData226-1 DData227-1 DData228-1 DData229-1 DData230-1 DData231-1 DData232-1 DData233-1 DData234-1 DData235-1 DData236-1 DData237-1 DData238-1 DData239-1 Data240-1 Data241-1 Data242-1 Data243-1 Data244-1 Data245-1 Data246-1 Data247-1 Data248-1 Data249-1 Data250-1 Data251-1 Data252-1 Data253-1 Data254-1 Data255-1 Out0-2-1 Out1-2-1 Out2-2-1 Out3-2-1 Out4-2-1 Out5-2-1 Out6-2-1 Out7-2-1 Out8-2-1	RoyalRoad

x35	Req1-2	Ready1-2	Fitness-Estimation-Ack-Pin1-2 DData0-2 DData1-2 DData2-2 DData3-2 DData4-2 DData5-2 DData6-2 DData7-2 DData8-2 DData9-2 DData10-2 DData11-2 DData12-2 DData13-2 DData14-2 DData15-2 Data16-2 Data17-2 Data18-2 Data19-2 Data20-2 Data21-2 Data22-2 Data23-2 Data24-2 Data25-2 Data26-2 Data27-2 Data28-2 Data29-2 Data30-2 Data31-2 DData32-2 DData33-2 DData34-2 DData35-2 DData36-2 DData37-2 DData38-2 DData39-2 DData40-2 DData41-2 DData42-2 DData43-2 DData44-2 DData45-2 DData46-2 DData47-2 Data48-2 Data49-2 Data50-2 Data51-2 Data52-2 Data53-2 Data54-2 Data55-2 Data56-2 Data57-2 Data58-2 Data59-2 Data60-2 Data61-2 Data62-2 Data63-2 DData64-2 DData65-2 DData66-2 DData67-2 DData68-2 DData69-2 DData70-2 DData71-2 DData72-2 DData73-2 DData74-2 DData75-2 DData76-2 DData77-2 DData78-2 DData79-2 Data80-2 Data81-2 Data82-2 Data83-2 Data84-2 Data85-2 Data86-2 Data87-2 Data88-2 Data89-2 Data90-2 Data91-2 Data92-2 Data93-2 Data94-2 Data95-2 DData96-2 DData97-2 DData98-2 DData99-2 DData100-2 DData101-2 DData102-2 DData103-2 DData104-2 DData105-2 DData106-2 DData107-2 DData108-2 DData109-2 DData110-2 DData111-2 Data112-2 Data113-2 Data114-2 Data115-2 Data116-2 Data117-2 Data118-2 Data119-2 Data120-2 Data121-2 Data122-2 Data123-2 Data124-2 Data125-2 Data126-2 Data127-2 DData128-2 DData129-2 DData130-2 DData131-2 DData132-2 DData133-2 DData134-2 DData135-2 DData136-2 DData137-2 DData138-2 DData139-2 DData140-2 DData141-2 DData142-2 DData143-2 Data144-2 Data145-2 Data146-2 Data147-2 Data148-2 Data149-2 Data150-2 Data151-2 Data152-2 Data153-2 Data154-2 Data155-2 Data156-2 Data157-2 Data158-2 Data159-2 DData160-2 DData161-2 DData162-2 DData163-2 DData164-2 DData165-2 DData166-2 DData167-2 DData168-2 DData169-2 DData170-2 DData171-2 DData172-2 DData173-2 DData174-2 DData175-2 Data176-2 Data177-2 Data178-2 Data179-2 Data180-2 Data181-2 Data182-2 Data183-2 Data184-2 Data185-2 Data186-2 Data187-2 Data188-2 Data189-2 Data190-2 Data191-2 DData192-2 DData193-2 DData194-2 DData195-2 DData196-2 DData197-2 DData198-2 DData199-2 DData200-2 DData201-2 DData202-2 DData203-2 DData204-2 DData205-2 DData206-2 DData207-2 Data208-2 Data209-2 Data210-2 Data211-2 Data212-2 Data213-2 Data214-2 Data215-2 Data216-2 Data217-2 Data218-2 Data219-2 Data220-2 Data221-2 Data222-2 Data223-2 DData224-2 DData225-2 DData226-2 DData227-2 DData228-2 DData229-2 DData230-2 DData231-2 DData232-2 DData233-2 DData234-2 DData235-2 DData236-2 DData237-2 DData238-2 DData239-2 Data240-2 Data241-2 Data242-2 Data243-2 Data244-2 Data245-2 Data246-2 Data247-2 Data248-2 Data249-2 Data250-2 Data251-2 Data252-2 Data253-2 Data254-2 Data255-2 Out0-1-2 Out1-1-2 Out2-1-2 Out3-1-2 Out4-1-2 Out5-1-2 Out6-1-2 Out7-1-2 Out8-1-2	RoyalRoad
x36	Req2-2	Ready2-2	Fitness-Estimation-Ack-Pin2-2 DData0-2 DData1-2 DData2-2 DData3-2 DData4-2 DData5-2 DData6-2 DData7-2 DData8-2 DData9-2 DData10-2 DData11-2 DData12-2 DData13-2 DData14-2 DData15-2 Data16-2 Data17-2 Data18-2 Data19-2 Data20-2 Data21-2 Data22-2 Data23-2 Data24-2 Data25-2 Data26-2 Data27-2 Data28-2 Data29-2 Data30-2 Data31-2 DData32-2 DData33-2 DData34-2 DData35-2 DData36-2 DData37-2 DData38-2 DData39-2 DData40-2 DData41-2 DData42-2 DData43-2 DData44-2 DData45-2 DData46-2 DData47-2 Data48-2 Data49-2 Data50-2 Data51-2 Data52-2 Data53-2 Data54-2 Data55-2 Data56-2 Data57-2 Data58-2 Data59-2 Data60-2 Data61-2 Data62-2 Data63-2 DData64-2 DData65-2 DData66-2 DData67-2 DData68-2 DData69-2 DData70-2 DData71-2 DData72-2 DData73-2 DData74-2 DData75-2 DData76-2 DData77-2 DData78-2 DData79-2 Data80-2 Data81-2 Data82-2 Data83-2 Data84-2 Data85-2 Data86-2 Data87-2 Data88-2 Data89-2 Data90-2 Data91-2 Data92-2 Data93-2 Data94-2 Data95-2 DData96-2 DData97-2 DData98-2 DData99-2 DData100-2 DData101-2 DData102-2 DData103-2 DData104-2 DData105-2 DData106-2 DData107-2 DData108-2 DData109-2 DData110-2 DData111-2 Data112-2 Data113-2 Data114-2 Data115-2 Data116-2 Data117-2 Data118-2 Data119-2 Data120-2 Data121-2 Data122-2 Data123-2 Data124-2 Data125-2 Data126-2 Data127-2 DData128-2 DData129-2 DData130-2 DData131-2 DData132-2 DData133-2 DData134-2 DData135-2 DData136-2 DData137-2 DData138-2 DData139-2 DData140-2 DData141-2 DData142-2 DData143-2 Data144-2 Data145-2 Data146-2 Data147-2 Data148-2 Data149-2 Data150-2 Data151-2 Data152-2 Data153-2 Data154-2 Data155-2 Data156-2 Data157-2 Data158-2 Data159-2 DData160-2 DData161-2 DData162-2 DData163-2 DData164-2 DData165-2 DData166-2 DData167-2 DData168-2 DData169-2 DData170-2 DData171-2 DData172-2 DData173-2 DData174-2 DData175-2 Data176-2 Data177-2 Data178-2 Data179-2 Data180-2 Data181-2 Data182-2 Data183-2 Data184-2 Data185-2 Data186-2 Data187-2 Data188-2 Data189-2 Data190-2 Data191-2 DData192-2 DData193-2 DData194-2 DData195-2 DData196-2 DData197-2 DData198-2 DData199-2 DData200-2 DData201-2 DData202-2 DData203-2 DData204-2 DData205-2 DData206-2 DData207-2 Data208-2 Data209-2 Data210-2 Data211-2 Data212-2 Data213-2 Data214-2 Data215-2 Data216-2 Data217-2 Data218-2 Data219-2 Data220-2 Data221-2 Data222-2 Data223-2 DData224-2 DData225-2 DData226-2 DData227-2 DData228-2 DData229-2 DData230-2 DData231-2 DData232-2 DData233-2 DData234-2 DData235-2 DData236-2 DData237-2 DData238-2 DData239-2 Data240-2 Data241-2 Data242-2 Data243-2 Data244-2 Data245-2 Data246-2 Data247-2 Data248-2 Data249-2 Data250-2 Data251-2 Data252-2 Data253-2 Data254-2 Data255-2 Out0-2-2 Out1-2-2 Out2-2-2 Out3-2-2 Out4-2-2 Out5-2-2 Out6-2-2 Out7-2-2 Out8-2-2	RoyalRoad

x37	Req1-3	Ready1-3	Fitness-Estimation-Ack-Pin1-3 DData0-3 DData1-3 DData2-3 DData3-3 DData4-3 DData5-3 DData6-3 DData7-3 DData8-3 DData9-3 DData10-3 DData11-3 DData12-3 DData13-3 DData14-3 DData15-3 Data16-3 Data17-3 Data18-3 Data19-3 Data20-3 Data21-3 Data22-3 Data23-3 Data24-3 Data25-3 Data26-3 Data27-3 Data28-3 Data29-3 Data30-3 Data31-3 DData32-3 DData33-3 DData34-3 DData35-3 DData36-3 DData37-3 DData38-3 DData39-3 DData40-3 DData41-3 DData42-3 DData43-3 DData44-3 DData45-3 DData46-3 DData47-3 Data48-3 Data49-3 Data50-3 Data51-3 Data52-3 Data53-3 Data54-3 Data55-3 Data56-3 Data57-3 Data58-3 Data59-3 Data60-3 Data61-3 Data62-3 Data63-3 DData64-3 DData65-3 DData66-3 DData67-3 DData68-3 DData69-3 DData70-3 DData71-3 DData72-3 DData73-3 DData74-3 DData75-3 DData76-3 DData77-3 DData78-3 DData79-3 Data80-3 Data81-3 Data82-3 Data83-3 Data84-3 Data85-3 Data86-3 Data87-3 Data88-3 Data89-3 Data90-3 Data91-3 Data92-3 Data93-3 Data94-3 Data95-3 DData96-3 DData97-3 DData98-3 DData99-3 DData100-3 DData101-3 DData102-3 DData103-3 DData104-3 DData105-3 DData106-3 DData107-3 DData108-3 DData109-3 DData110-3 DData111-3 Data112-3 Data113-3 Data114-3 Data115-3 Data116-3 Data117-3 Data118-3 Data119-3 Data120-3 Data121-3 Data122-3 Data123-3 Data124-3 Data125-3 Data126-3 Data127-3 DData128-3 DData129-3 DData130-3 DData131-3 DData132-3 DData133-3 DData134-3 DData135-3 DData136-3 DData137-3 DData138-3 DData139-3 DData140-3 DData141-3 DData142-3 DData143-3 Data144-3 Data145-3 Data146-3 Data147-3 Data148-3 Data149-3 Data150-3 Data151-3 Data152-3 Data153-3 Data154-3 Data155-3 Data156-3 Data157-3 Data158-3 Data159-3 DData160-3 DData161-3 DData162-3 DData163-3 DData164-3 DData165-3 DData166-3 DData167-3 DData168-3 DData169-3 DData170-3 DData171-3 DData172-3 DData173-3 DData174-3 DData175-3 Data176-3 Data177-3 Data178-3 Data179-3 Data180-3 Data181-3 Data182-3 Data183-3 Data184-3 Data185-3 Data186-3 Data187-3 Data188-3 Data189-3 Data190-3 Data191-3 DData192-3 DData193-3 DData194-3 DData195-3 DData196-3 DData197-3 DData198-3 DData199-3 DData200-3 DData201-3 DData202-3 DData203-3 DData204-3 DData205-3 DData206-3 DData207-3 Data208-3 Data209-3 Data210-3 Data211-3 Data212-3 Data213-3 Data214-3 Data215-3 Data216-3 Data217-3 Data218-3 Data219-3 Data220-3 Data221-3 Data222-3 Data223-3 DData224-3 DData225-3 DData226-3 DData227-3 DData228-3 DData229-3 DData230-3 DData231-3 DData232-3 DData233-3 DData234-3 DData235-3 DData236-3 DData237-3 DData238-3 DData239-3 Data240-3 Data241-3 Data242-3 Data243-3 Data244-3 Data245-3 Data246-3 Data247-3 Data248-3 Data249-3 Data250-3 Data251-3 Data252-3 Data253-3 Data254-3 Data255-3 Out0-1-3 Out1-1-3 Out2-1-3 Out3-1-3 Out4-1-3 Out5-1-3 Out6-1-3 Out7-1-3 Out8-1-3	RoyalRoad
x38	Req2-3	Ready2-3	Fitness-Estimation-Ack-Pin2-3 DData0-3 DData1-3 DData2-3 DData3-3 DData4-3 DData5-3 DData6-3 DData7-3 DData8-3 DData9-3 DData10-3 DData11-3 DData12-3 DData13-3 DData14-3 DData15-3 Data16-3 Data17-3 Data18-3 Data19-3 Data20-3 Data21-3 Data22-3 Data23-3 Data24-3 Data25-3 Data26-3 Data27-3 Data28-3 Data29-3 Data30-3 Data31-3 DData32-3 DData33-3 DData34-3 DData35-3 DData36-3 DData37-3 DData38-3 DData39-3 DData40-3 DData41-3 DData42-3 DData43-3 DData44-3 DData45-3 DData46-3 DData47-3 Data48-3 Data49-3 Data50-3 Data51-3 Data52-3 Data53-3 Data54-3 Data55-3 Data56-3 Data57-3 Data58-3 Data59-3 Data60-3 Data61-3 Data62-3 Data63-3 DData64-3 DData65-3 DData66-3 DData67-3 DData68-3 DData69-3 DData70-3 DData71-3 DData72-3 DData73-3 DData74-3 DData75-3 DData76-3 DData77-3 DData78-3 DData79-3 Data80-3 Data81-3 Data82-3 Data83-3 Data84-3 Data85-3 Data86-3 Data87-3 Data88-3 Data89-3 Data90-3 Data91-3 Data92-3 Data93-3 Data94-3 Data95-3 DData96-3 DData97-3 DData98-3 DData99-3 DData100-3 DData101-3 DData102-3 DData103-3 DData104-3 DData105-3 DData106-3 DData107-3 DData108-3 DData109-3 DData110-3 DData111-3 Data112-3 Data113-3 Data114-3 Data115-3 Data116-3 Data117-3 Data118-3 Data119-3 Data120-3 Data121-3 Data122-3 Data123-3 Data124-3 Data125-3 Data126-3 Data127-3 DData128-3 DData129-3 DData130-3 DData131-3 DData132-3 DData133-3 DData134-3 DData135-3 DData136-3 DData137-3 DData138-3 DData139-3 DData140-3 DData141-3 DData142-3 DData143-3 Data144-3 Data145-3 Data146-3 Data147-3 Data148-3 Data149-3 Data150-3 Data151-3 Data152-3 Data153-3 Data154-3 Data155-3 Data156-3 Data157-3 Data158-3 Data159-3 DData160-3 DData161-3 DData162-3 DData163-3 DData164-3 DData165-3 DData166-3 DData167-3 DData168-3 DData169-3 DData170-3 DData171-3 DData172-3 DData173-3 DData174-3 DData175-3 Data176-3 Data177-3 Data178-3 Data179-3 Data180-3 Data181-3 Data182-3 Data183-3 Data184-3 Data185-3 Data186-3 Data187-3 Data188-3 Data189-3 Data190-3 Data191-3 DData192-3 DData193-3 DData194-3 DData195-3 DData196-3 DData197-3 DData198-3 DData199-3 DData200-3 DData201-3 DData202-3 DData203-3 DData204-3 DData205-3 DData206-3 DData207-3 Data208-3 Data209-3 Data210-3 Data211-3 Data212-3 Data213-3 Data214-3 Data215-3 Data216-3 Data217-3 Data218-3 Data219-3 Data220-3 Data221-3 Data222-3 Data223-3 DData224-3 DData225-3 DData226-3 DData227-3 DData228-3 DData229-3 DData230-3 DData231-3 DData232-3 DData233-3 DData234-3 DData235-3 DData236-3 DData237-3 DData238-3 DData239-3 Data240-3 Data241-3 Data242-3 Data243-3 Data244-3 Data245-3 Data246-3 Data247-3 Data248-3 Data249-3 Data250-3 Data251-3 Data252-3 Data253-3 Data254-3 Data255-3 Out0-2-3 Out1-2-3 Out2-2-3 Out3-2-3 Out4-2-3 Out5-2-3 Out6-2-3 Out7-2-3 Out8-2-3	RoyalRoad

x39	Req1-4	Ready1-4	Fitness-Estimation-Ack-Pin1-4 DData0-4 DData1-4 DData2-4 DData3-4 DData4-4 DData5-4 DData6-4 DData7-4 DData8-4 DData9-4 DData10-4 DData11-4 DData12-4 DData13-4 DData14-4 DData15-4 Data16-4 Data17-4 Data18-4 Data19-4 Data20-4 Data21-4 Data22-4 Data23-4 Data24-4 Data25-4 Data26-4 Data27-4 Data28-4 Data29-4 Data30-4 Data31-4 DData32-4 DData33-4 DData34-4 DData35-4 DData36-4 DData37-4 DData38-4 DData39-4 DData40-4 DData41-4 DData42-4 DData43-4 DData44-4 DData45-4 DData46-4 DData47-4 Data48-4 Data49-4 Data50-4 Data51-4 Data52-4 Data53-4 Data54-4 Data55-4 Data56-4 Data57-4 Data58-4 Data59-4 Data60-4 Data61-4 Data62-4 Data63-4 DData64-4 DData65-4 DData66-4 DData67-4 DData68-4 DData69-4 DData70-4 DData71-4 DData72-4 DData73-4 DData74-4 DData75-4 DData76-4 DData77-4 DData78-4 DData79-4 Data80-4 Data81-4 Data82-4 Data83-4 Data84-4 Data85-4 Data86-4 Data87-4 Data88-4 Data89-4 Data90-4 Data91-4 Data92-4 Data93-4 Data94-4 Data95-4 DData96-4 DData97-4 DData98-4 DData99-4 DData100-4 DData101-4 DData102-4 DData103-4 DData104-4 DData105-4 DData106-4 DData107-4 DData108-4 DData109-4 DData110-4 DData111-4 Data112-4 Data113-4 Data114-4 Data115-4 Data116-4 Data117-4 Data118-4 Data119-4 Data120-4 Data121-4 Data122-4 Data123-4 Data124-4 Data125-4 Data126-4 Data127-4 DData128-4 DData129-4 DData130-4 DData131-4 DData132-4 DData133-4 DData134-4 DData135-4 DData136-4 DData137-4 DData138-4 DData139-4 DData140-4 DData141-4 DData142-4 DData143-4 Data144-4 Data145-4 Data146-4 Data147-4 Data148-4 Data149-4 Data150-4 Data151-4 Data152-4 Data153-4 Data154-4 Data155-4 Data156-4 Data157-4 Data158-4 Data159-4 DData160-4 DData161-4 DData162-4 DData163-4 DData164-4 DData165-4 DData166-4 DData167-4 DData168-4 DData169-4 DData170-4 DData171-4 DData172-4 DData173-4 DData174-4 DData175-4 Data176-4 Data177-4 Data178-4 Data179-4 Data180-4 Data181-4 Data182-4 Data183-4 Data184-4 Data185-4 Data186-4 Data187-4 Data188-4 Data189-4 Data190-4 Data191-4 DData192-4 DData193-4 DData194-4 DData195-4 DData196-4 DData197-4 DData198-4 DData199-4 DData200-4 DData201-4 DData202-4 DData203-4 DData204-4 DData205-4 DData206-4 DData207-4 Data208-4 Data209-4 Data210-4 Data211-4 Data212-4 Data213-4 Data214-4 Data215-4 Data216-4 Data217-4 Data218-4 Data219-4 Data220-4 Data221-4 Data222-4 Data223-4 DData224-4 DData225-4 DData226-4 DData227-4 DData228-4 DData229-4 DData230-4 DData231-4 DData232-4 DData233-4 DData234-4 DData235-4 DData236-4 DData237-4 DData238-4 DData239-4 Data240-4 Data241-4 Data242-4 Data243-4 Data244-4 Data245-4 Data246-4 Data247-4 Data248-4 Data249-4 Data250-4 Data251-4 Data252-4 Data253-4 Data254-4 Data255-4 Out0-1-4 Out1-1-4 Out2-1-4 Out3-1-4 Out4-1-4 Out5-1-4 Out6-1-4 Out7-1-4 Out8-1-4	RoyalRoad
x40	Req2-4	Ready2-4	Fitness-Estimation-Ack-Pin2-4 DData0-4 DData1-4 DData2-4 DData3-4 DData4-4 DData5-4 DData6-4 DData7-4 DData8-4 DData9-4 DData10-4 DData11-4 DData12-4 DData13-4 DData14-4 DData15-4 Data16-4 Data17-4 Data18-4 Data19-4 Data20-4 Data21-4 Data22-4 Data23-4 Data24-4 Data25-4 Data26-4 Data27-4 Data28-4 Data29-4 Data30-4 Data31-4 DData32-4 DData33-4 DData34-4 DData35-4 DData36-4 DData37-4 DData38-4 DData39-4 DData40-4 DData41-4 DData42-4 DData43-4 DData44-4 DData45-4 DData46-4 DData47-4 Data48-4 Data49-4 Data50-4 Data51-4 Data52-4 Data53-4 Data54-4 Data55-4 Data56-4 Data57-4 Data58-4 Data59-4 Data60-4 Data61-4 Data62-4 Data63-4 DData64-4 DData65-4 DData66-4 DData67-4 DData68-4 DData69-4 DData70-4 DData71-4 DData72-4 DData73-4 DData74-4 DData75-4 DData76-4 DData77-4 DData78-4 DData79-4 Data80-4 Data81-4 Data82-4 Data83-4 Data84-4 Data85-4 Data86-4 Data87-4 Data88-4 Data89-4 Data90-4 Data91-4 Data92-4 Data93-4 Data94-4 Data95-4 DData96-4 DData97-4 DData98-4 DData99-4 DData100-4 DData101-4 DData102-4 DData103-4 DData104-4 DData105-4 DData106-4 DData107-4 DData108-4 DData109-4 DData110-4 DData111-4 Data112-4 Data113-4 Data114-4 Data115-4 Data116-4 Data117-4 Data118-4 Data119-4 Data120-4 Data121-4 Data122-4 Data123-4 Data124-4 Data125-4 Data126-4 Data127-4 DData128-4 DData129-4 DData130-4 DData131-4 DData132-4 DData133-4 DData134-4 DData135-4 DData136-4 DData137-4 DData138-4 DData139-4 DData140-4 DData141-4 DData142-4 DData143-4 Data144-4 Data145-4 Data146-4 Data147-4 Data148-4 Data149-4 Data150-4 Data151-4 Data152-4 Data153-4 Data154-4 Data155-4 Data156-4 Data157-4 Data158-4 Data159-4 DData160-4 DData161-4 DData162-4 DData163-4 DData164-4 DData165-4 DData166-4 DData167-4 DData168-4 DData169-4 DData170-4 DData171-4 DData172-4 DData173-4 DData174-4 DData175-4 Data176-4 Data177-4 Data178-4 Data179-4 Data180-4 Data181-4 Data182-4 Data183-4 Data184-4 Data185-4 Data186-4 Data187-4 Data188-4 Data189-4 Data190-4 Data191-4 DData192-4 DData193-4 DData194-4 DData195-4 DData196-4 DData197-4 DData198-4 DData199-4 DData200-4 DData201-4 DData202-4 DData203-4 DData204-4 DData205-4 DData206-4 DData207-4 Data208-4 Data209-4 Data210-4 Data211-4 Data212-4 Data213-4 Data214-4 Data215-4 Data216-4 Data217-4 Data218-4 Data219-4 Data220-4 Data221-4 Data222-4 Data223-4 DData224-4 DData225-4 DData226-4 DData227-4 DData228-4 DData229-4 DData230-4 DData231-4 DData232-4 DData233-4 DData234-4 DData235-4 DData236-4 DData237-4 DData238-4 DData239-4 Data240-4 Data241-4 Data242-4 Data243-4 Data244-4 Data245-4 Data246-4 Data247-4 Data248-4 Data249-4 Data250-4 Data251-4 Data252-4 Data253-4 Data254-4 Data255-4 Out0-2-4 Out1-2-4 Out2-2-4 Out3-2-4 Out4-2-4 Out5-2-4 Out6-2-4 Out7-2-4 Out8-2-4	RoyalRoad


******External Circuit
**Fitness Function I/O Data Bus Switch
x41	out0-1-1 out1-1-1 out2-1-1 out3-1-1 out4-1-1 out5-1-1 out6-1-1 out7-1-1 out8-1-1 0 0 0 0 0 0 0 	out0-1-1 out1-1-1 out2-1-1 out3-1-1 out4-1-1 out5-1-1 out6-1-1 out7-1-1 out8-1-1 0 0 0 0 0 0 0 	out0-1-1 out1-1-1 out2-1-1 out3-1-1 out4-1-1 out5-1-1 out6-1-1 out7-1-1 out8-1-1 0 0 0 0 0 0 0 	out0-1-1 out1-1-1 out2-1-1 out3-1-1 out4-1-1 out5-1-1 out6-1-1 out7-1-1 out8-1-1 0 0 0 0 0 0 0 	out0-1-1 out1-1-1 out2-1-1 out3-1-1 out4-1-1 out5-1-1 out6-1-1 out7-1-1 out8-1-1 0 0 0 0 0 0 0 	out0-1-1 out1-1-1 out2-1-1 out3-1-1 out4-1-1 out5-1-1 out6-1-1 out7-1-1 out8-1-1 0 0 0 0 0 0 0 	out0-1-1 out1-1-1 out2-1-1 out3-1-1 out4-1-1 out5-1-1 out6-1-1 out7-1-1 out8-1-1 0 0 0 0 0 0 0 	out0-1-1 out1-1-1 out2-1-1 out3-1-1 out4-1-1 out5-1-1 out6-1-1 out7-1-1 out8-1-1 0 0 0 0 0 0 0 	DData0-1 DData1-1 DData2-1 DData3-1 DData4-1 DData5-1 DData6-1 DData7-1 DData8-1 DData9-1 DData10-1 DData11-1 DData12-1 DData13-1 DData14-1 DData15-1 DData32-1 DData33-1 DData34-1 DData35-1 DData36-1 DData37-1 DData38-1 DData39-1 DData40-1 DData41-1 DData42-1 DData43-1 DData44-1 DData45-1 DData46-1 DData47-1 DData64-1 DData65-1 DData66-1 DData67-1 DData68-1 DData69-1 DData70-1 DData71-1 DData72-1 DData73-1 DData74-1 DData75-1 DData76-1 DData77-1 DData78-1 DData79-1 DData96-1 DData97-1 DData98-1 DData99-1 DData100-1 DData101-1 DData102-1 DData103-1 DData104-1 DData105-1 DData106-1 DData107-1 DData108-1 DData109-1 DData110-1 DData111-1 DData128-1 DData129-1 DData130-1 DData131-1 DData132-1 DData133-1 DData134-1 DData135-1 DData136-1 DData137-1 DData138-1 DData139-1 DData140-1 DData141-1 DData142-1 DData143-1 DData160-1 DData161-1 DData162-1 DData163-1 DData164-1 DData165-1 DData166-1 DData167-1 DData168-1 DData169-1 DData170-1 DData171-1 DData172-1 DData173-1 DData174-1 DData175-1 DData192-1 DData193-1 DData194-1 DData195-1 DData196-1 DData197-1 DData198-1 DData199-1 DData200-1 DData201-1 DData202-1 DData203-1 DData204-1 DData205-1 DData206-1 DData207-1 DData224-1 DData225-1 DData226-1 DData227-1 DData228-1 DData229-1 DData230-1 DData231-1 DData232-1 DData233-1 DData234-1 DData235-1 DData236-1 DData237-1 DData238-1 DData239-1	preData0-1 preData1-1 preData2-1 preData3-1 preData4-1 preData5-1 preData6-1 preData7-1 preData8-1 preData9-1 preData10-1 preData11-1 preData12-1 preData13-1 preData14-1 preData15-1 preData16-1 preData17-1 preData18-1 preData19-1 preData20-1 preData21-1 preData22-1 preData23-1 preData24-1 preData25-1 preData26-1 preData27-1 preData28-1 preData29-1 preData30-1 preData31-1 preData32-1 preData33-1 preData34-1 preData35-1 preData36-1 preData37-1 preData38-1 preData39-1 preData40-1 preData41-1 preData42-1 preData43-1 preData44-1 preData45-1 preData46-1 preData47-1 preData48-1 preData49-1 preData50-1 preData51-1 preData52-1 preData53-1 preData54-1 preData55-1 preData56-1 preData57-1 preData58-1 preData59-1 preData60-1 preData61-1 preData62-1 preData63-1 preData64-1 preData65-1 preData66-1 preData67-1 preData68-1 preData69-1 preData70-1 preData71-1 preData72-1 preData73-1 preData74-1 preData75-1 preData76-1 preData77-1 preData78-1 preData79-1 preData80-1 preData81-1 preData82-1 preData83-1 preData84-1 preData85-1 preData86-1 preData87-1 preData88-1 preData89-1 preData90-1 preData91-1 preData92-1 preData93-1 preData94-1 preData95-1 preData96-1 preData97-1 preData98-1 preData99-1 preData100-1 preData101-1 preData102-1 preData103-1 preData104-1 preData105-1 preData106-1 preData107-1 preData108-1 preData109-1 preData110-1 preData111-1 preData112-1 preData113-1 preData114-1 preData115-1 preData116-1 preData117-1 preData118-1 preData119-1 preData120-1 preData121-1 preData122-1 preData123-1 preData124-1 preData125-1 preData126-1 preData127-1	Ready1-1	Ready1-1^	MUX-Array-128-no-INV	wn=3u	wp=9u	*m=20
x42	out0-2-1 out1-2-1 out2-2-1 out3-2-1 out4-2-1 out5-2-1 out6-2-1 out7-2-1 out8-2-1 0 0 0 0 0 0 0 	out0-2-1 out1-2-1 out2-2-1 out3-2-1 out4-2-1 out5-2-1 out6-2-1 out7-2-1 out8-2-1 0 0 0 0 0 0 0 	out0-2-1 out1-2-1 out2-2-1 out3-2-1 out4-2-1 out5-2-1 out6-2-1 out7-2-1 out8-2-1 0 0 0 0 0 0 0 	out0-2-1 out1-2-1 out2-2-1 out3-2-1 out4-2-1 out5-2-1 out6-2-1 out7-2-1 out8-2-1 0 0 0 0 0 0 0 	out0-2-1 out1-2-1 out2-2-1 out3-2-1 out4-2-1 out5-2-1 out6-2-1 out7-2-1 out8-2-1 0 0 0 0 0 0 0 	out0-2-1 out1-2-1 out2-2-1 out3-2-1 out4-2-1 out5-2-1 out6-2-1 out7-2-1 out8-2-1 0 0 0 0 0 0 0 	out0-2-1 out1-2-1 out2-2-1 out3-2-1 out4-2-1 out5-2-1 out6-2-1 out7-2-1 out8-2-1 0 0 0 0 0 0 0 	out0-2-1 out1-2-1 out2-2-1 out3-2-1 out4-2-1 out5-2-1 out6-2-1 out7-2-1 out8-2-1 0 0 0 0 0 0 0 	preData0-1 preData1-1 preData2-1 preData3-1 preData4-1 preData5-1 preData6-1 preData7-1 preData8-1 preData9-1 preData10-1 preData11-1 preData12-1 preData13-1 preData14-1 preData15-1 preData16-1 preData17-1 preData18-1 preData19-1 preData20-1 preData21-1 preData22-1 preData23-1 preData24-1 preData25-1 preData26-1 preData27-1 preData28-1 preData29-1 preData30-1 preData31-1 preData32-1 preData33-1 preData34-1 preData35-1 preData36-1 preData37-1 preData38-1 preData39-1 preData40-1 preData41-1 preData42-1 preData43-1 preData44-1 preData45-1 preData46-1 preData47-1 preData48-1 preData49-1 preData50-1 preData51-1 preData52-1 preData53-1 preData54-1 preData55-1 preData56-1 preData57-1 preData58-1 preData59-1 preData60-1 preData61-1 preData62-1 preData63-1 preData64-1 preData65-1 preData66-1 preData67-1 preData68-1 preData69-1 preData70-1 preData71-1 preData72-1 preData73-1 preData74-1 preData75-1 preData76-1 preData77-1 preData78-1 preData79-1 preData80-1 preData81-1 preData82-1 preData83-1 preData84-1 preData85-1 preData86-1 preData87-1 preData88-1 preData89-1 preData90-1 preData91-1 preData92-1 preData93-1 preData94-1 preData95-1 preData96-1 preData97-1 preData98-1 preData99-1 preData100-1 preData101-1 preData102-1 preData103-1 preData104-1 preData105-1 preData106-1 preData107-1 preData108-1 preData109-1 preData110-1 preData111-1 preData112-1 preData113-1 preData114-1 preData115-1 preData116-1 preData117-1 preData118-1 preData119-1 preData120-1 preData121-1 preData122-1 preData123-1 preData124-1 preData125-1 preData126-1 preData127-1	Data0-1 Data1-1 Data2-1 Data3-1 Data4-1 Data5-1 Data6-1 Data7-1 Data8-1 Data9-1 Data10-1 Data11-1 Data12-1 Data13-1 Data14-1 Data15-1 Data32-1 Data33-1 Data34-1 Data35-1 Data36-1 Data37-1 Data38-1 Data39-1 Data40-1 Data41-1 Data42-1 Data43-1 Data44-1 Data45-1 Data46-1 Data47-1 Data64-1 Data65-1 Data66-1 Data67-1 Data68-1 Data69-1 Data70-1 Data71-1 Data72-1 Data73-1 Data74-1 Data75-1 Data76-1 Data77-1 Data78-1 Data79-1 Data96-1 Data97-1 Data98-1 Data99-1 Data100-1 Data101-1 Data102-1 Data103-1 Data104-1 Data105-1 Data106-1 Data107-1 Data108-1 Data109-1 Data110-1 Data111-1 Data128-1 Data129-1 Data130-1 Data131-1 Data132-1 Data133-1 Data134-1 Data135-1 Data136-1 Data137-1 Data138-1 Data139-1 Data140-1 Data141-1 Data142-1 Data143-1 Data160-1 Data161-1 Data162-1 Data163-1 Data164-1 Data165-1 Data166-1 Data167-1 Data168-1 Data169-1 Data170-1 Data171-1 Data172-1 Data173-1 Data174-1 Data175-1 Data192-1 Data193-1 Data194-1 Data195-1 Data196-1 Data197-1 Data198-1 Data199-1 Data200-1 Data201-1 Data202-1 Data203-1 Data204-1 Data205-1 Data206-1 Data207-1 Data224-1 Data225-1 Data226-1 Data227-1 Data228-1 Data229-1 Data230-1 Data231-1 Data232-1 Data233-1 Data234-1 Data235-1 Data236-1 Data237-1 Data238-1 Data239-1	Ready2-1	Ready2-1^	MUX-Array-128-no-INV	wn=3u	wp=9u	*m=20

x43	out0-1-2 out1-1-2 out2-1-2 out3-1-2 out4-1-2 out5-1-2 out6-1-2 out7-1-2 out8-1-2 0 0 0 0 0 0 0 	out0-1-2 out1-1-2 out2-1-2 out3-1-2 out4-1-2 out5-1-2 out6-1-2 out7-1-2 out8-1-2 0 0 0 0 0 0 0 	out0-1-2 out1-1-2 out2-1-2 out3-1-2 out4-1-2 out5-1-2 out6-1-2 out7-1-2 out8-1-2 0 0 0 0 0 0 0 	out0-1-2 out1-1-2 out2-1-2 out3-1-2 out4-1-2 out5-1-2 out6-1-2 out7-1-2 out8-1-2 0 0 0 0 0 0 0 	out0-1-2 out1-1-2 out2-1-2 out3-1-2 out4-1-2 out5-1-2 out6-1-2 out7-1-2 out8-1-2 0 0 0 0 0 0 0 	out0-1-2 out1-1-2 out2-1-2 out3-1-2 out4-1-2 out5-1-2 out6-1-2 out7-1-2 out8-1-2 0 0 0 0 0 0 0 	out0-1-2 out1-1-2 out2-1-2 out3-1-2 out4-1-2 out5-1-2 out6-1-2 out7-1-2 out8-1-2 0 0 0 0 0 0 0 	out0-1-2 out1-1-2 out2-1-2 out3-1-2 out4-1-2 out5-1-2 out6-1-2 out7-1-2 out8-1-2 0 0 0 0 0 0 0 	DData0-2 DData1-2 DData2-2 DData3-2 DData4-2 DData5-2 DData6-2 DData7-2 DData8-2 DData9-2 DData10-2 DData11-2 DData12-2 DData13-2 DData14-2 DData15-2 DData32-2 DData33-2 DData34-2 DData35-2 DData36-2 DData37-2 DData38-2 DData39-2 DData40-2 DData41-2 DData42-2 DData43-2 DData44-2 DData45-2 DData46-2 DData47-2 DData64-2 DData65-2 DData66-2 DData67-2 DData68-2 DData69-2 DData70-2 DData71-2 DData72-2 DData73-2 DData74-2 DData75-2 DData76-2 DData77-2 DData78-2 DData79-2 DData96-2 DData97-2 DData98-2 DData99-2 DData100-2 DData101-2 DData102-2 DData103-2 DData104-2 DData105-2 DData106-2 DData107-2 DData108-2 DData109-2 DData110-2 DData111-2 DData128-2 DData129-2 DData130-2 DData131-2 DData132-2 DData133-2 DData134-2 DData135-2 DData136-2 DData137-2 DData138-2 DData139-2 DData140-2 DData141-2 DData142-2 DData143-2 DData160-2 DData161-2 DData162-2 DData163-2 DData164-2 DData165-2 DData166-2 DData167-2 DData168-2 DData169-2 DData170-2 DData171-2 DData172-2 DData173-2 DData174-2 DData175-2 DData192-2 DData193-2 DData194-2 DData195-2 DData196-2 DData197-2 DData198-2 DData199-2 DData200-2 DData201-2 DData202-2 DData203-2 DData204-2 DData205-2 DData206-2 DData207-2 DData224-2 DData225-2 DData226-2 DData227-2 DData228-2 DData229-2 DData230-2 DData231-2 DData232-2 DData233-2 DData234-2 DData235-2 DData236-2 DData237-2 DData238-2 DData239-2	preData0-2 preData1-2 preData2-2 preData3-2 preData4-2 preData5-2 preData6-2 preData7-2 preData8-2 preData9-2 preData10-2 preData11-2 preData12-2 preData13-2 preData14-2 preData15-2 preData16-2 preData17-2 preData18-2 preData19-2 preData20-2 preData21-2 preData22-2 preData23-2 preData24-2 preData25-2 preData26-2 preData27-2 preData28-2 preData29-2 preData30-2 preData31-2 preData32-2 preData33-2 preData34-2 preData35-2 preData36-2 preData37-2 preData38-2 preData39-2 preData40-2 preData41-2 preData42-2 preData43-2 preData44-2 preData45-2 preData46-2 preData47-2 preData48-2 preData49-2 preData50-2 preData51-2 preData52-2 preData53-2 preData54-2 preData55-2 preData56-2 preData57-2 preData58-2 preData59-2 preData60-2 preData61-2 preData62-2 preData63-2 preData64-2 preData65-2 preData66-2 preData67-2 preData68-2 preData69-2 preData70-2 preData71-2 preData72-2 preData73-2 preData74-2 preData75-2 preData76-2 preData77-2 preData78-2 preData79-2 preData80-2 preData81-2 preData82-2 preData83-2 preData84-2 preData85-2 preData86-2 preData87-2 preData88-2 preData89-2 preData90-2 preData91-2 preData92-2 preData93-2 preData94-2 preData95-2 preData96-2 preData97-2 preData98-2 preData99-2 preData100-2 preData101-2 preData102-2 preData103-2 preData104-2 preData105-2 preData106-2 preData107-2 preData108-2 preData109-2 preData110-2 preData111-2 preData112-2 preData113-2 preData114-2 preData115-2 preData116-2 preData117-2 preData118-2 preData119-2 preData120-2 preData121-2 preData122-2 preData123-2 preData124-2 preData125-2 preData126-2 preData127-2	Ready1-2	Ready1-2^	MUX-Array-128-no-INV	wn=3u	wp=9u	*m=20
x44	out0-2-2 out1-2-2 out2-2-2 out3-2-2 out4-2-2 out5-2-2 out6-2-2 out7-2-2 out8-2-2 0 0 0 0 0 0 0 	out0-2-2 out1-2-2 out2-2-2 out3-2-2 out4-2-2 out5-2-2 out6-2-2 out7-2-2 out8-2-2 0 0 0 0 0 0 0 	out0-2-2 out1-2-2 out2-2-2 out3-2-2 out4-2-2 out5-2-2 out6-2-2 out7-2-2 out8-2-2 0 0 0 0 0 0 0 	out0-2-2 out1-2-2 out2-2-2 out3-2-2 out4-2-2 out5-2-2 out6-2-2 out7-2-2 out8-2-2 0 0 0 0 0 0 0 	out0-2-2 out1-2-2 out2-2-2 out3-2-2 out4-2-2 out5-2-2 out6-2-2 out7-2-2 out8-2-2 0 0 0 0 0 0 0 	out0-2-2 out1-2-2 out2-2-2 out3-2-2 out4-2-2 out5-2-2 out6-2-2 out7-2-2 out8-2-2 0 0 0 0 0 0 0 	out0-2-2 out1-2-2 out2-2-2 out3-2-2 out4-2-2 out5-2-2 out6-2-2 out7-2-2 out8-2-2 0 0 0 0 0 0 0 	out0-2-2 out1-2-2 out2-2-2 out3-2-2 out4-2-2 out5-2-2 out6-2-2 out7-2-2 out8-2-2 0 0 0 0 0 0 0 	preData0-2 preData1-2 preData2-2 preData3-2 preData4-2 preData5-2 preData6-2 preData7-2 preData8-2 preData9-2 preData10-2 preData11-2 preData12-2 preData13-2 preData14-2 preData15-2 preData16-2 preData17-2 preData18-2 preData19-2 preData20-2 preData21-2 preData22-2 preData23-2 preData24-2 preData25-2 preData26-2 preData27-2 preData28-2 preData29-2 preData30-2 preData31-2 preData32-2 preData33-2 preData34-2 preData35-2 preData36-2 preData37-2 preData38-2 preData39-2 preData40-2 preData41-2 preData42-2 preData43-2 preData44-2 preData45-2 preData46-2 preData47-2 preData48-2 preData49-2 preData50-2 preData51-2 preData52-2 preData53-2 preData54-2 preData55-2 preData56-2 preData57-2 preData58-2 preData59-2 preData60-2 preData61-2 preData62-2 preData63-2 preData64-2 preData65-2 preData66-2 preData67-2 preData68-2 preData69-2 preData70-2 preData71-2 preData72-2 preData73-2 preData74-2 preData75-2 preData76-2 preData77-2 preData78-2 preData79-2 preData80-2 preData81-2 preData82-2 preData83-2 preData84-2 preData85-2 preData86-2 preData87-2 preData88-2 preData89-2 preData90-2 preData91-2 preData92-2 preData93-2 preData94-2 preData95-2 preData96-2 preData97-2 preData98-2 preData99-2 preData100-2 preData101-2 preData102-2 preData103-2 preData104-2 preData105-2 preData106-2 preData107-2 preData108-2 preData109-2 preData110-2 preData111-2 preData112-2 preData113-2 preData114-2 preData115-2 preData116-2 preData117-2 preData118-2 preData119-2 preData120-2 preData121-2 preData122-2 preData123-2 preData124-2 preData125-2 preData126-2 preData127-2	Data0-2 Data1-2 Data2-2 Data3-2 Data4-2 Data5-2 Data6-2 Data7-2 Data8-2 Data9-2 Data10-2 Data11-2 Data12-2 Data13-2 Data14-2 Data15-2 Data32-2 Data33-2 Data34-2 Data35-2 Data36-2 Data37-2 Data38-2 Data39-2 Data40-2 Data41-2 Data42-2 Data43-2 Data44-2 Data45-2 Data46-2 Data47-2 Data64-2 Data65-2 Data66-2 Data67-2 Data68-2 Data69-2 Data70-2 Data71-2 Data72-2 Data73-2 Data74-2 Data75-2 Data76-2 Data77-2 Data78-2 Data79-2 Data96-2 Data97-2 Data98-2 Data99-2 Data100-2 Data101-2 Data102-2 Data103-2 Data104-2 Data105-2 Data106-2 Data107-2 Data108-2 Data109-2 Data110-2 Data111-2 Data128-2 Data129-2 Data130-2 Data131-2 Data132-2 Data133-2 Data134-2 Data135-2 Data136-2 Data137-2 Data138-2 Data139-2 Data140-2 Data141-2 Data142-2 Data143-2 Data160-2 Data161-2 Data162-2 Data163-2 Data164-2 Data165-2 Data166-2 Data167-2 Data168-2 Data169-2 Data170-2 Data171-2 Data172-2 Data173-2 Data174-2 Data175-2 Data192-2 Data193-2 Data194-2 Data195-2 Data196-2 Data197-2 Data198-2 Data199-2 Data200-2 Data201-2 Data202-2 Data203-2 Data204-2 Data205-2 Data206-2 Data207-2 Data224-2 Data225-2 Data226-2 Data227-2 Data228-2 Data229-2 Data230-2 Data231-2 Data232-2 Data233-2 Data234-2 Data235-2 Data236-2 Data237-2 Data238-2 Data239-2	Ready2-2	Ready2-2^	MUX-Array-128-no-INV	wn=3u	wp=9u	*m=20

x45	out0-1-3 out1-1-3 out2-1-3 out3-1-3 out4-1-3 out5-1-3 out6-1-3 out7-1-3 out8-1-3 0 0 0 0 0 0 0 	out0-1-3 out1-1-3 out2-1-3 out3-1-3 out4-1-3 out5-1-3 out6-1-3 out7-1-3 out8-1-3 0 0 0 0 0 0 0 	out0-1-3 out1-1-3 out2-1-3 out3-1-3 out4-1-3 out5-1-3 out6-1-3 out7-1-3 out8-1-3 0 0 0 0 0 0 0 	out0-1-3 out1-1-3 out2-1-3 out3-1-3 out4-1-3 out5-1-3 out6-1-3 out7-1-3 out8-1-3 0 0 0 0 0 0 0 	out0-1-3 out1-1-3 out2-1-3 out3-1-3 out4-1-3 out5-1-3 out6-1-3 out7-1-3 out8-1-3 0 0 0 0 0 0 0 	out0-1-3 out1-1-3 out2-1-3 out3-1-3 out4-1-3 out5-1-3 out6-1-3 out7-1-3 out8-1-3 0 0 0 0 0 0 0 	out0-1-3 out1-1-3 out2-1-3 out3-1-3 out4-1-3 out5-1-3 out6-1-3 out7-1-3 out8-1-3 0 0 0 0 0 0 0 	out0-1-3 out1-1-3 out2-1-3 out3-1-3 out4-1-3 out5-1-3 out6-1-3 out7-1-3 out8-1-3 0 0 0 0 0 0 0 	DData0-3 DData1-3 DData2-3 DData3-3 DData4-3 DData5-3 DData6-3 DData7-3 DData8-3 DData9-3 DData10-3 DData11-3 DData12-3 DData13-3 DData14-3 DData15-3 DData32-3 DData33-3 DData34-3 DData35-3 DData36-3 DData37-3 DData38-3 DData39-3 DData40-3 DData41-3 DData42-3 DData43-3 DData44-3 DData45-3 DData46-3 DData47-3 DData64-3 DData65-3 DData66-3 DData67-3 DData68-3 DData69-3 DData70-3 DData71-3 DData72-3 DData73-3 DData74-3 DData75-3 DData76-3 DData77-3 DData78-3 DData79-3 DData96-3 DData97-3 DData98-3 DData99-3 DData100-3 DData101-3 DData102-3 DData103-3 DData104-3 DData105-3 DData106-3 DData107-3 DData108-3 DData109-3 DData110-3 DData111-3 DData128-3 DData129-3 DData130-3 DData131-3 DData132-3 DData133-3 DData134-3 DData135-3 DData136-3 DData137-3 DData138-3 DData139-3 DData140-3 DData141-3 DData142-3 DData143-3 DData160-3 DData161-3 DData162-3 DData163-3 DData164-3 DData165-3 DData166-3 DData167-3 DData168-3 DData169-3 DData170-3 DData171-3 DData172-3 DData173-3 DData174-3 DData175-3 DData192-3 DData193-3 DData194-3 DData195-3 DData196-3 DData197-3 DData198-3 DData199-3 DData200-3 DData201-3 DData202-3 DData203-3 DData204-3 DData205-3 DData206-3 DData207-3 DData224-3 DData225-3 DData226-3 DData227-3 DData228-3 DData229-3 DData230-3 DData231-3 DData232-3 DData233-3 DData234-3 DData235-3 DData236-3 DData237-3 DData238-3 DData239-3	preData0-3 preData1-3 preData2-3 preData3-3 preData4-3 preData5-3 preData6-3 preData7-3 preData8-3 preData9-3 preData10-3 preData11-3 preData12-3 preData13-3 preData14-3 preData15-3 preData16-3 preData17-3 preData18-3 preData19-3 preData20-3 preData21-3 preData22-3 preData23-3 preData24-3 preData25-3 preData26-3 preData27-3 preData28-3 preData29-3 preData30-3 preData31-3 preData32-3 preData33-3 preData34-3 preData35-3 preData36-3 preData37-3 preData38-3 preData39-3 preData40-3 preData41-3 preData42-3 preData43-3 preData44-3 preData45-3 preData46-3 preData47-3 preData48-3 preData49-3 preData50-3 preData51-3 preData52-3 preData53-3 preData54-3 preData55-3 preData56-3 preData57-3 preData58-3 preData59-3 preData60-3 preData61-3 preData62-3 preData63-3 preData64-3 preData65-3 preData66-3 preData67-3 preData68-3 preData69-3 preData70-3 preData71-3 preData72-3 preData73-3 preData74-3 preData75-3 preData76-3 preData77-3 preData78-3 preData79-3 preData80-3 preData81-3 preData82-3 preData83-3 preData84-3 preData85-3 preData86-3 preData87-3 preData88-3 preData89-3 preData90-3 preData91-3 preData92-3 preData93-3 preData94-3 preData95-3 preData96-3 preData97-3 preData98-3 preData99-3 preData100-3 preData101-3 preData102-3 preData103-3 preData104-3 preData105-3 preData106-3 preData107-3 preData108-3 preData109-3 preData110-3 preData111-3 preData112-3 preData113-3 preData114-3 preData115-3 preData116-3 preData117-3 preData118-3 preData119-3 preData120-3 preData121-3 preData122-3 preData123-3 preData124-3 preData125-3 preData126-3 preData127-3	Ready1-3	Ready1-3^	MUX-Array-128-no-INV	wn=3u	wp=9u	*m=20
x46	out0-2-3 out1-2-3 out2-2-3 out3-2-3 out4-2-3 out5-2-3 out6-2-3 out7-2-3 out8-2-3 0 0 0 0 0 0 0 	out0-2-3 out1-2-3 out2-2-3 out3-2-3 out4-2-3 out5-2-3 out6-2-3 out7-2-3 out8-2-3 0 0 0 0 0 0 0 	out0-2-3 out1-2-3 out2-2-3 out3-2-3 out4-2-3 out5-2-3 out6-2-3 out7-2-3 out8-2-3 0 0 0 0 0 0 0 	out0-2-3 out1-2-3 out2-2-3 out3-2-3 out4-2-3 out5-2-3 out6-2-3 out7-2-3 out8-2-3 0 0 0 0 0 0 0 	out0-2-3 out1-2-3 out2-2-3 out3-2-3 out4-2-3 out5-2-3 out6-2-3 out7-2-3 out8-2-3 0 0 0 0 0 0 0 	out0-2-3 out1-2-3 out2-2-3 out3-2-3 out4-2-3 out5-2-3 out6-2-3 out7-2-3 out8-2-3 0 0 0 0 0 0 0 	out0-2-3 out1-2-3 out2-2-3 out3-2-3 out4-2-3 out5-2-3 out6-2-3 out7-2-3 out8-2-3 0 0 0 0 0 0 0 	out0-2-3 out1-2-3 out2-2-3 out3-2-3 out4-2-3 out5-2-3 out6-2-3 out7-2-3 out8-2-3 0 0 0 0 0 0 0 	preData0-3 preData1-3 preData2-3 preData3-3 preData4-3 preData5-3 preData6-3 preData7-3 preData8-3 preData9-3 preData10-3 preData11-3 preData12-3 preData13-3 preData14-3 preData15-3 preData16-3 preData17-3 preData18-3 preData19-3 preData20-3 preData21-3 preData22-3 preData23-3 preData24-3 preData25-3 preData26-3 preData27-3 preData28-3 preData29-3 preData30-3 preData31-3 preData32-3 preData33-3 preData34-3 preData35-3 preData36-3 preData37-3 preData38-3 preData39-3 preData40-3 preData41-3 preData42-3 preData43-3 preData44-3 preData45-3 preData46-3 preData47-3 preData48-3 preData49-3 preData50-3 preData51-3 preData52-3 preData53-3 preData54-3 preData55-3 preData56-3 preData57-3 preData58-3 preData59-3 preData60-3 preData61-3 preData62-3 preData63-3 preData64-3 preData65-3 preData66-3 preData67-3 preData68-3 preData69-3 preData70-3 preData71-3 preData72-3 preData73-3 preData74-3 preData75-3 preData76-3 preData77-3 preData78-3 preData79-3 preData80-3 preData81-3 preData82-3 preData83-3 preData84-3 preData85-3 preData86-3 preData87-3 preData88-3 preData89-3 preData90-3 preData91-3 preData92-3 preData93-3 preData94-3 preData95-3 preData96-3 preData97-3 preData98-3 preData99-3 preData100-3 preData101-3 preData102-3 preData103-3 preData104-3 preData105-3 preData106-3 preData107-3 preData108-3 preData109-3 preData110-3 preData111-3 preData112-3 preData113-3 preData114-3 preData115-3 preData116-3 preData117-3 preData118-3 preData119-3 preData120-3 preData121-3 preData122-3 preData123-3 preData124-3 preData125-3 preData126-3 preData127-3	Data0-3 Data1-3 Data2-3 Data3-3 Data4-3 Data5-3 Data6-3 Data7-3 Data8-3 Data9-3 Data10-3 Data11-3 Data12-3 Data13-3 Data14-3 Data15-3 Data32-3 Data33-3 Data34-3 Data35-3 Data36-3 Data37-3 Data38-3 Data39-3 Data40-3 Data41-3 Data42-3 Data43-3 Data44-3 Data45-3 Data46-3 Data47-3 Data64-3 Data65-3 Data66-3 Data67-3 Data68-3 Data69-3 Data70-3 Data71-3 Data72-3 Data73-3 Data74-3 Data75-3 Data76-3 Data77-3 Data78-3 Data79-3 Data96-3 Data97-3 Data98-3 Data99-3 Data100-3 Data101-3 Data102-3 Data103-3 Data104-3 Data105-3 Data106-3 Data107-3 Data108-3 Data109-3 Data110-3 Data111-3 Data128-3 Data129-3 Data130-3 Data131-3 Data132-3 Data133-3 Data134-3 Data135-3 Data136-3 Data137-3 Data138-3 Data139-3 Data140-3 Data141-3 Data142-3 Data143-3 Data160-3 Data161-3 Data162-3 Data163-3 Data164-3 Data165-3 Data166-3 Data167-3 Data168-3 Data169-3 Data170-3 Data171-3 Data172-3 Data173-3 Data174-3 Data175-3 Data192-3 Data193-3 Data194-3 Data195-3 Data196-3 Data197-3 Data198-3 Data199-3 Data200-3 Data201-3 Data202-3 Data203-3 Data204-3 Data205-3 Data206-3 Data207-3 Data224-3 Data225-3 Data226-3 Data227-3 Data228-3 Data229-3 Data230-3 Data231-3 Data232-3 Data233-3 Data234-3 Data235-3 Data236-3 Data237-3 Data238-3 Data239-3	Ready2-3	Ready2-3^	MUX-Array-128-no-INV	wn=3u	wp=9u	*m=20

x47	out0-1-4 out1-1-4 out2-1-4 out3-1-4 out4-1-4 out5-1-4 out6-1-4 out7-1-4 out8-1-4 0 0 0 0 0 0 0 	out0-1-4 out1-1-4 out2-1-4 out3-1-4 out4-1-4 out5-1-4 out6-1-4 out7-1-4 out8-1-4 0 0 0 0 0 0 0 	out0-1-4 out1-1-4 out2-1-4 out3-1-4 out4-1-4 out5-1-4 out6-1-4 out7-1-4 out8-1-4 0 0 0 0 0 0 0 	out0-1-4 out1-1-4 out2-1-4 out3-1-4 out4-1-4 out5-1-4 out6-1-4 out7-1-4 out8-1-4 0 0 0 0 0 0 0 	out0-1-4 out1-1-4 out2-1-4 out3-1-4 out4-1-4 out5-1-4 out6-1-4 out7-1-4 out8-1-4 0 0 0 0 0 0 0 	out0-1-4 out1-1-4 out2-1-4 out3-1-4 out4-1-4 out5-1-4 out6-1-4 out7-1-4 out8-1-4 0 0 0 0 0 0 0 	out0-1-4 out1-1-4 out2-1-4 out3-1-4 out4-1-4 out5-1-4 out6-1-4 out7-1-4 out8-1-4 0 0 0 0 0 0 0 	out0-1-4 out1-1-4 out2-1-4 out3-1-4 out4-1-4 out5-1-4 out6-1-4 out7-1-4 out8-1-4 0 0 0 0 0 0 0 	DData0-4 DData1-4 DData2-4 DData3-4 DData4-4 DData5-4 DData6-4 DData7-4 DData8-4 DData9-4 DData10-4 DData11-4 DData12-4 DData13-4 DData14-4 DData15-4 DData32-4 DData33-4 DData34-4 DData35-4 DData36-4 DData37-4 DData38-4 DData39-4 DData40-4 DData41-4 DData42-4 DData43-4 DData44-4 DData45-4 DData46-4 DData47-4 DData64-4 DData65-4 DData66-4 DData67-4 DData68-4 DData69-4 DData70-4 DData71-4 DData72-4 DData73-4 DData74-4 DData75-4 DData76-4 DData77-4 DData78-4 DData79-4 DData96-4 DData97-4 DData98-4 DData99-4 DData100-4 DData101-4 DData102-4 DData103-4 DData104-4 DData105-4 DData106-4 DData107-4 DData108-4 DData109-4 DData110-4 DData111-4 DData128-4 DData129-4 DData130-4 DData131-4 DData132-4 DData133-4 DData134-4 DData135-4 DData136-4 DData137-4 DData138-4 DData139-4 DData140-4 DData141-4 DData142-4 DData143-4 DData160-4 DData161-4 DData162-4 DData163-4 DData164-4 DData165-4 DData166-4 DData167-4 DData168-4 DData169-4 DData170-4 DData171-4 DData172-4 DData173-4 DData174-4 DData175-4 DData192-4 DData193-4 DData194-4 DData195-4 DData196-4 DData197-4 DData198-4 DData199-4 DData200-4 DData201-4 DData202-4 DData203-4 DData204-4 DData205-4 DData206-4 DData207-4 DData224-4 DData225-4 DData226-4 DData227-4 DData228-4 DData229-4 DData230-4 DData231-4 DData232-4 DData233-4 DData234-4 DData235-4 DData236-4 DData237-4 DData238-4 DData239-4	preData0-4 preData1-4 preData2-4 preData3-4 preData4-4 preData5-4 preData6-4 preData7-4 preData8-4 preData9-4 preData10-4 preData11-4 preData12-4 preData13-4 preData14-4 preData15-4 preData16-4 preData17-4 preData18-4 preData19-4 preData20-4 preData21-4 preData22-4 preData23-4 preData24-4 preData25-4 preData26-4 preData27-4 preData28-4 preData29-4 preData30-4 preData31-4 preData32-4 preData33-4 preData34-4 preData35-4 preData36-4 preData37-4 preData38-4 preData39-4 preData40-4 preData41-4 preData42-4 preData43-4 preData44-4 preData45-4 preData46-4 preData47-4 preData48-4 preData49-4 preData50-4 preData51-4 preData52-4 preData53-4 preData54-4 preData55-4 preData56-4 preData57-4 preData58-4 preData59-4 preData60-4 preData61-4 preData62-4 preData63-4 preData64-4 preData65-4 preData66-4 preData67-4 preData68-4 preData69-4 preData70-4 preData71-4 preData72-4 preData73-4 preData74-4 preData75-4 preData76-4 preData77-4 preData78-4 preData79-4 preData80-4 preData81-4 preData82-4 preData83-4 preData84-4 preData85-4 preData86-4 preData87-4 preData88-4 preData89-4 preData90-4 preData91-4 preData92-4 preData93-4 preData94-4 preData95-4 preData96-4 preData97-4 preData98-4 preData99-4 preData100-4 preData101-4 preData102-4 preData103-4 preData104-4 preData105-4 preData106-4 preData107-4 preData108-4 preData109-4 preData110-4 preData111-4 preData112-4 preData113-4 preData114-4 preData115-4 preData116-4 preData117-4 preData118-4 preData119-4 preData120-4 preData121-4 preData122-4 preData123-4 preData124-4 preData125-4 preData126-4 preData127-4	Ready1-4	Ready1-4^	MUX-Array-128-no-INV	wn=3u	wp=9u	*m=20
x48	out0-2-4 out1-2-4 out2-2-4 out3-2-4 out4-2-4 out5-2-4 out6-2-4 out7-2-4 out8-2-4 0 0 0 0 0 0 0 	out0-2-4 out1-2-4 out2-2-4 out3-2-4 out4-2-4 out5-2-4 out6-2-4 out7-2-4 out8-2-4 0 0 0 0 0 0 0 	out0-2-4 out1-2-4 out2-2-4 out3-2-4 out4-2-4 out5-2-4 out6-2-4 out7-2-4 out8-2-4 0 0 0 0 0 0 0 	out0-2-4 out1-2-4 out2-2-4 out3-2-4 out4-2-4 out5-2-4 out6-2-4 out7-2-4 out8-2-4 0 0 0 0 0 0 0 	out0-2-4 out1-2-4 out2-2-4 out3-2-4 out4-2-4 out5-2-4 out6-2-4 out7-2-4 out8-2-4 0 0 0 0 0 0 0 	out0-2-4 out1-2-4 out2-2-4 out3-2-4 out4-2-4 out5-2-4 out6-2-4 out7-2-4 out8-2-4 0 0 0 0 0 0 0 	out0-2-4 out1-2-4 out2-2-4 out3-2-4 out4-2-4 out5-2-4 out6-2-4 out7-2-4 out8-2-4 0 0 0 0 0 0 0 	out0-2-4 out1-2-4 out2-2-4 out3-2-4 out4-2-4 out5-2-4 out6-2-4 out7-2-4 out8-2-4 0 0 0 0 0 0 0 	preData0-4 preData1-4 preData2-4 preData3-4 preData4-4 preData5-4 preData6-4 preData7-4 preData8-4 preData9-4 preData10-4 preData11-4 preData12-4 preData13-4 preData14-4 preData15-4 preData16-4 preData17-4 preData18-4 preData19-4 preData20-4 preData21-4 preData22-4 preData23-4 preData24-4 preData25-4 preData26-4 preData27-4 preData28-4 preData29-4 preData30-4 preData31-4 preData32-4 preData33-4 preData34-4 preData35-4 preData36-4 preData37-4 preData38-4 preData39-4 preData40-4 preData41-4 preData42-4 preData43-4 preData44-4 preData45-4 preData46-4 preData47-4 preData48-4 preData49-4 preData50-4 preData51-4 preData52-4 preData53-4 preData54-4 preData55-4 preData56-4 preData57-4 preData58-4 preData59-4 preData60-4 preData61-4 preData62-4 preData63-4 preData64-4 preData65-4 preData66-4 preData67-4 preData68-4 preData69-4 preData70-4 preData71-4 preData72-4 preData73-4 preData74-4 preData75-4 preData76-4 preData77-4 preData78-4 preData79-4 preData80-4 preData81-4 preData82-4 preData83-4 preData84-4 preData85-4 preData86-4 preData87-4 preData88-4 preData89-4 preData90-4 preData91-4 preData92-4 preData93-4 preData94-4 preData95-4 preData96-4 preData97-4 preData98-4 preData99-4 preData100-4 preData101-4 preData102-4 preData103-4 preData104-4 preData105-4 preData106-4 preData107-4 preData108-4 preData109-4 preData110-4 preData111-4 preData112-4 preData113-4 preData114-4 preData115-4 preData116-4 preData117-4 preData118-4 preData119-4 preData120-4 preData121-4 preData122-4 preData123-4 preData124-4 preData125-4 preData126-4 preData127-4	Data0-4 Data1-4 Data2-4 Data3-4 Data4-4 Data5-4 Data6-4 Data7-4 Data8-4 Data9-4 Data10-4 Data11-4 Data12-4 Data13-4 Data14-4 Data15-4 Data32-4 Data33-4 Data34-4 Data35-4 Data36-4 Data37-4 Data38-4 Data39-4 Data40-4 Data41-4 Data42-4 Data43-4 Data44-4 Data45-4 Data46-4 Data47-4 Data64-4 Data65-4 Data66-4 Data67-4 Data68-4 Data69-4 Data70-4 Data71-4 Data72-4 Data73-4 Data74-4 Data75-4 Data76-4 Data77-4 Data78-4 Data79-4 Data96-4 Data97-4 Data98-4 Data99-4 Data100-4 Data101-4 Data102-4 Data103-4 Data104-4 Data105-4 Data106-4 Data107-4 Data108-4 Data109-4 Data110-4 Data111-4 Data128-4 Data129-4 Data130-4 Data131-4 Data132-4 Data133-4 Data134-4 Data135-4 Data136-4 Data137-4 Data138-4 Data139-4 Data140-4 Data141-4 Data142-4 Data143-4 Data160-4 Data161-4 Data162-4 Data163-4 Data164-4 Data165-4 Data166-4 Data167-4 Data168-4 Data169-4 Data170-4 Data171-4 Data172-4 Data173-4 Data174-4 Data175-4 Data192-4 Data193-4 Data194-4 Data195-4 Data196-4 Data197-4 Data198-4 Data199-4 Data200-4 Data201-4 Data202-4 Data203-4 Data204-4 Data205-4 Data206-4 Data207-4 Data224-4 Data225-4 Data226-4 Data227-4 Data228-4 Data229-4 Data230-4 Data231-4 Data232-4 Data233-4 Data234-4 Data235-4 Data236-4 Data237-4 Data238-4 Data239-4	Ready2-4	Ready2-4^	MUX-Array-128-no-INV	wn=3u	wp=9u	*m=20


*AND Gates for Req. and Ready Signals
x49	Fitness-Estimation-Ready1-Pad1-1	Fitness-Estimation-Ready1-Pad2-1	Fitness-Estimation-Ready1-Pad3-1	Fitness-Estimation-Ready1-Pad4-1	Fitness-Estimation-Ready1-Pad5-1	Fitness-Estimation-Ready1-Pad6-1	Fitness-Estimation-Ready1-Pad7-1	Fitness-Estimation-Ready1-Pad8-1	Ready1-1	Ready1-1^	AND8-m20	wn=16u	wp=48u	*m=20
x50	Fitness-Estimation-Ready2-Pad1-1	Fitness-Estimation-Ready2-Pad2-1	Fitness-Estimation-Ready2-Pad3-1	Fitness-Estimation-Ready2-Pad4-1	Fitness-Estimation-Ready2-Pad5-1	Fitness-Estimation-Ready2-Pad6-1	Fitness-Estimation-Ready2-Pad7-1	Fitness-Estimation-Ready2-Pad8-1	Ready2-1	Ready2-1^	AND8-m20	wn=16u	wp=48u	*m=20
x51	Fitness-Estimation-Req1-Pad1-1	Fitness-Estimation-Req1-Pad2-1	Fitness-Estimation-Req1-Pad3-1	Fitness-Estimation-Req1-Pad4-1	Fitness-Estimation-Req1-Pad5-1	Fitness-Estimation-Req1-Pad6-1	Fitness-Estimation-Req1-Pad7-1	Fitness-Estimation-Req1-Pad8-1	Req1-1	Req1-1^	AND8-m20	wn=16u	wp=48u	*m=20
x52	Fitness-Estimation-Req2-Pad1-1	Fitness-Estimation-Req2-Pad2-1	Fitness-Estimation-Req2-Pad3-1	Fitness-Estimation-Req2-Pad4-1	Fitness-Estimation-Req2-Pad5-1	Fitness-Estimation-Req2-Pad6-1	Fitness-Estimation-Req2-Pad7-1	Fitness-Estimation-Req2-Pad8-1	Req2-1	Req2-1^	AND8-m20	wn=16u	wp=48u	*m=20

x53	Fitness-Estimation-Ready1-Pad1-2	Fitness-Estimation-Ready1-Pad2-2	Fitness-Estimation-Ready1-Pad3-2	Fitness-Estimation-Ready1-Pad4-2	Fitness-Estimation-Ready1-Pad5-2	Fitness-Estimation-Ready1-Pad6-2	Fitness-Estimation-Ready1-Pad7-2	Fitness-Estimation-Ready1-Pad8-2	Ready1-2	Ready1-2^	AND8-m20	wn=16u	wp=48u	*m=20
x54	Fitness-Estimation-Ready2-Pad1-2	Fitness-Estimation-Ready2-Pad2-2	Fitness-Estimation-Ready2-Pad3-2	Fitness-Estimation-Ready2-Pad4-2	Fitness-Estimation-Ready2-Pad5-2	Fitness-Estimation-Ready2-Pad6-2	Fitness-Estimation-Ready2-Pad7-2	Fitness-Estimation-Ready2-Pad8-2	Ready2-2	Ready2-2^	AND8-m20	wn=16u	wp=48u	*m=20
x55	Fitness-Estimation-Req1-Pad1-2	Fitness-Estimation-Req1-Pad2-2	Fitness-Estimation-Req1-Pad3-2	Fitness-Estimation-Req1-Pad4-2	Fitness-Estimation-Req1-Pad5-2	Fitness-Estimation-Req1-Pad6-2	Fitness-Estimation-Req1-Pad7-2	Fitness-Estimation-Req1-Pad8-2	Req1-2	Req1-2^	AND8-m20	wn=16u	wp=48u	*m=20
x56	Fitness-Estimation-Req2-Pad1-2	Fitness-Estimation-Req2-Pad2-2	Fitness-Estimation-Req2-Pad3-2	Fitness-Estimation-Req2-Pad4-2	Fitness-Estimation-Req2-Pad5-2	Fitness-Estimation-Req2-Pad6-2	Fitness-Estimation-Req2-Pad7-2	Fitness-Estimation-Req2-Pad8-2	Req2-2	Req2-2^	AND8-m20	wn=16u	wp=48u	*m=20

x57	Fitness-Estimation-Ready1-Pad1-3	Fitness-Estimation-Ready1-Pad2-3	Fitness-Estimation-Ready1-Pad3-3	Fitness-Estimation-Ready1-Pad4-3	Fitness-Estimation-Ready1-Pad5-3	Fitness-Estimation-Ready1-Pad6-3	Fitness-Estimation-Ready1-Pad7-3	Fitness-Estimation-Ready1-Pad8-3	Ready1-3	Ready1-3^	AND8-m20	wn=16u	wp=48u	*m=20
x58	Fitness-Estimation-Ready2-Pad1-3	Fitness-Estimation-Ready2-Pad2-3	Fitness-Estimation-Ready2-Pad3-3	Fitness-Estimation-Ready2-Pad4-3	Fitness-Estimation-Ready2-Pad5-3	Fitness-Estimation-Ready2-Pad6-3	Fitness-Estimation-Ready2-Pad7-3	Fitness-Estimation-Ready2-Pad8-3	Ready2-3	Ready2-3^	AND8-m20	wn=16u	wp=48u	*m=20
x59	Fitness-Estimation-Req1-Pad1-3	Fitness-Estimation-Req1-Pad2-3	Fitness-Estimation-Req1-Pad3-3	Fitness-Estimation-Req1-Pad4-3	Fitness-Estimation-Req1-Pad5-3	Fitness-Estimation-Req1-Pad6-3	Fitness-Estimation-Req1-Pad7-3	Fitness-Estimation-Req1-Pad8-3	Req1-3	Req1-3^	AND8-m20	wn=16u	wp=48u	*m=20
x60	Fitness-Estimation-Req2-Pad1-3	Fitness-Estimation-Req2-Pad2-3	Fitness-Estimation-Req2-Pad3-3	Fitness-Estimation-Req2-Pad4-3	Fitness-Estimation-Req2-Pad5-3	Fitness-Estimation-Req2-Pad6-3	Fitness-Estimation-Req2-Pad7-3	Fitness-Estimation-Req2-Pad8-3	Req2-3	Req2-3^	AND8-m20	wn=16u	wp=48u	*m=20

x61	Fitness-Estimation-Ready1-Pad1-4	Fitness-Estimation-Ready1-Pad2-4	Fitness-Estimation-Ready1-Pad3-4	Fitness-Estimation-Ready1-Pad4-4	Fitness-Estimation-Ready1-Pad5-4	Fitness-Estimation-Ready1-Pad6-4	Fitness-Estimation-Ready1-Pad7-4	Fitness-Estimation-Ready1-Pad8-4	Ready1-4	Ready1-4^	AND8-m20	wn=16u	wp=48u	*m=20
x62	Fitness-Estimation-Ready2-Pad1-4	Fitness-Estimation-Ready2-Pad2-4	Fitness-Estimation-Ready2-Pad3-4	Fitness-Estimation-Ready2-Pad4-4	Fitness-Estimation-Ready2-Pad5-4	Fitness-Estimation-Ready2-Pad6-4	Fitness-Estimation-Ready2-Pad7-4	Fitness-Estimation-Ready2-Pad8-4	Ready2-4	Ready2-4^	AND8-m20	wn=16u	wp=48u	*m=20
x63	Fitness-Estimation-Req1-Pad1-4	Fitness-Estimation-Req1-Pad2-4	Fitness-Estimation-Req1-Pad3-4	Fitness-Estimation-Req1-Pad4-4	Fitness-Estimation-Req1-Pad5-4	Fitness-Estimation-Req1-Pad6-4	Fitness-Estimation-Req1-Pad7-4	Fitness-Estimation-Req1-Pad8-4	Req1-4	Req1-4^	AND8-m20	wn=16u	wp=48u	*m=20
x64	Fitness-Estimation-Req2-Pad1-4	Fitness-Estimation-Req2-Pad2-4	Fitness-Estimation-Req2-Pad3-4	Fitness-Estimation-Req2-Pad4-4	Fitness-Estimation-Req2-Pad5-4	Fitness-Estimation-Req2-Pad6-4	Fitness-Estimation-Req2-Pad7-4	Fitness-Estimation-Req2-Pad8-4	Req2-4	Req2-4^	AND8-m20	wn=16u	wp=48u	*m=20


*OR Gates for Fitness Unit Ack. Pins
x65	Fitness-Estimation-Ack-Pin1-1	Fitness-Estimation-Ack-Pin2-1	Fitness-Estimation-Ack-Pin-1	Fitness-Estimation-Ack-Pin-1^	OR2-m20	wn=16u	wp=48u	*m=20
x66	Fitness-Estimation-Ack-Pin1-2	Fitness-Estimation-Ack-Pin2-2	Fitness-Estimation-Ack-Pin-2	Fitness-Estimation-Ack-Pin-2^	OR2-m20	wn=16u	wp=48u	*m=20
x67	Fitness-Estimation-Ack-Pin1-3	Fitness-Estimation-Ack-Pin2-3	Fitness-Estimation-Ack-Pin-3	Fitness-Estimation-Ack-Pin-3^	OR2-m20	wn=16u	wp=48u	*m=20
x68	Fitness-Estimation-Ack-Pin1-4	Fitness-Estimation-Ack-Pin2-4	Fitness-Estimation-Ack-Pin-4	Fitness-Estimation-Ack-Pin-4^	OR2-m20	wn=16u	wp=48u	*m=20


*AND Gates for Multi-GAP Selection
x69	Selection-Ack-Pin2-1	Selection-Ack-Pin3-1	Selection-Ack-Pin4-1	Selection-Ack-Pin5-1	Selection-Ack-Pin6-1	Selection-Ack-Pin7-1	Selection-Ack-Pin8-1	vdd	Selection-Ack-Pin1-1	Selection-Ack-Pin1-1^	AND8-m20	wn=16u	wp=48u	*m=20	*Added a VDD input to use AND8 subcircuit for AND7
x70	Selection-Ack-Pin2-2	Selection-Ack-Pin3-2	Selection-Ack-Pin4-2	Selection-Ack-Pin5-2	Selection-Ack-Pin6-2	Selection-Ack-Pin7-2	Selection-Ack-Pin8-2	vdd	Selection-Ack-Pin1-2	Selection-Ack-Pin1-2^	AND8-m20	wn=16u	wp=48u	*m=20
x71	Selection-Ack-Pin2-3	Selection-Ack-Pin3-3	Selection-Ack-Pin4-3	Selection-Ack-Pin5-3	Selection-Ack-Pin6-3	Selection-Ack-Pin7-3	Selection-Ack-Pin8-3	vdd	Selection-Ack-Pin1-3	Selection-Ack-Pin1-3^	AND8-m20	wn=16u	wp=48u	*m=20
x72	Selection-Ack-Pin2-4	Selection-Ack-Pin3-4	Selection-Ack-Pin4-4	Selection-Ack-Pin5-4	Selection-Ack-Pin6-4	Selection-Ack-Pin7-4	Selection-Ack-Pin8-4	vdd	Selection-Ack-Pin1-4	Selection-Ack-Pin1-4^	AND8-m20	wn=16u	wp=48u	*m=20


******Components
***Array of 128 inverter-less multiplexers***
.subckt MUX-Array-128-no-INV	in0-1 in1-1 in2-1 in3-1 in4-1 in5-1 in6-1 in7-1 in8-1 in9-1 in10-1 in11-1 in12-1 in13-1 in14-1 in15-1 in16-1 in17-1 in18-1 in19-1 in20-1 in21-1 in22-1 in23-1 in24-1 in25-1 in26-1 in27-1 in28-1 in29-1 in30-1 in31-1 in32-1 in33-1 in34-1 in35-1 in36-1 in37-1 in38-1 in39-1 in40-1 in41-1 in42-1 in43-1 in44-1 in45-1 in46-1 in47-1 in48-1 in49-1 in50-1 in51-1 in52-1 in53-1 in54-1 in55-1 in56-1 in57-1 in58-1 in59-1 in60-1 in61-1 in62-1 in63-1 in64-1 in65-1 in66-1 in67-1 in68-1 in69-1 in70-1 in71-1 in72-1 in73-1 in74-1 in75-1 in76-1 in77-1 in78-1 in79-1 in80-1 in81-1 in82-1 in83-1 in84-1 in85-1 in86-1 in87-1 in88-1 in89-1 in90-1 in91-1 in92-1 in93-1 in94-1 in95-1 in96-1 in97-1 in98-1 in99-1 in100-1 in101-1 in102-1 in103-1 in104-1 in105-1 in106-1 in107-1 in108-1 in109-1 in110-1 in111-1 in112-1 in113-1 in114-1 in115-1 in116-1 in117-1 in118-1 in119-1 in120-1 in121-1 in122-1 in123-1 in124-1 in125-1 in126-1 in127-1	in0-2 in1-2 in2-2 in3-2 in4-2 in5-2 in6-2 in7-2 in8-2 in9-2 in10-2 in11-2 in12-2 in13-2 in14-2 in15-2 in16-2 in17-2 in18-2 in19-2 in20-2 in21-2 in22-2 in23-2 in24-2 in25-2 in26-2 in27-2 in28-2 in29-2 in30-2 in31-2 in32-2 in33-2 in34-2 in35-2 in36-2 in37-2 in38-2 in39-2 in40-2 in41-2 in42-2 in43-2 in44-2 in45-2 in46-2 in47-2 in48-2 in49-2 in50-2 in51-2 in52-2 in53-2 in54-2 in55-2 in56-2 in57-2 in58-2 in59-2 in60-2 in61-2 in62-2 in63-2 in64-2 in65-2 in66-2 in67-2 in68-2 in69-2 in70-2 in71-2 in72-2 in73-2 in74-2 in75-2 in76-2 in77-2 in78-2 in79-2 in80-2 in81-2 in82-2 in83-2 in84-2 in85-2 in86-2 in87-2 in88-2 in89-2 in90-2 in91-2 in92-2 in93-2 in94-2 in95-2 in96-2 in97-2 in98-2 in99-2 in100-2 in101-2 in102-2 in103-2 in104-2 in105-2 in106-2 in107-2 in108-2 in109-2 in110-2 in111-2 in112-2 in113-2 in114-2 in115-2 in116-2 in117-2 in118-2 in119-2 in120-2 in121-2 in122-2 in123-2 in124-2 in125-2 in126-2 in127-2	out0 out1 out2 out3 out4 out5 out6 out7 out8 out9 out10 out11 out12 out13 out14 out15 out16 out17 out18 out19 out20 out21 out22 out23 out24 out25 out26 out27 out28 out29 out30 out31 out32 out33 out34 out35 out36 out37 out38 out39 out40 out41 out42 out43 out44 out45 out46 out47 out48 out49 out50 out51 out52 out53 out54 out55 out56 out57 out58 out59 out60 out61 out62 out63 out64 out65 out66 out67 out68 out69 out70 out71 out72 out73 out74 out75 out76 out77 out78 out79 out80 out81 out82 out83 out84 out85 out86 out87 out88 out89 out90 out91 out92 out93 out94 out95 out96 out97 out98 out99 out100 out101 out102 out103 out104 out105 out106 out107 out108 out109 out110 out111 out112 out113 out114 out115 out116 out117 out118 out119 out120 out121 out122 out123 out124 out125 out126 out127	control	control^	wn=1u	wp=3u	le=0.18u
x1	in0-1 in1-1 in2-1 in3-1 in4-1 in5-1 in6-1 in7-1 in8-1 in9-1 in10-1 in11-1 in12-1 in13-1 in14-1 in15-1 in0-2 in1-2 in2-2 in3-2 in4-2 in5-2 in6-2 in7-2 in8-2 in9-2 in10-2 in11-2 in12-2 in13-2 in14-2 in15-2 out0 out1 out2 out3 out4 out5 out6 out7 out8 out9 out10 out11 out12 out13 out14 out15	control	control^	MUX-Array-16-no-INV	wn='wn'	wp='wp'	le='le'
x2	in16-1 in17-1 in18-1 in19-1 in20-1 in21-1 in22-1 in23-1 in24-1 in25-1 in26-1 in27-1 in28-1 in29-1 in30-1 in31-1 in16-2 in17-2 in18-2 in19-2 in20-2 in21-2 in22-2 in23-2 in24-2 in25-2 in26-2 in27-2 in28-2 in29-2 in30-2 in31-2 out16 out17 out18 out19 out20 out21 out22 out23 out24 out25 out26 out27 out28 out29 out30 out31	control	control^	MUX-Array-16-no-INV	wn='wn'	wp='wp'	le='le'
x3	in32-1 in33-1 in34-1 in35-1 in36-1 in37-1 in38-1 in39-1 in40-1 in41-1 in42-1 in43-1 in44-1 in45-1 in46-1 in47-1 in32-2 in33-2 in34-2 in35-2 in36-2 in37-2 in38-2 in39-2 in40-2 in41-2 in42-2 in43-2 in44-2 in45-2 in46-2 in47-2 out32 out33 out34 out35 out36 out37 out38 out39 out40 out41 out42 out43 out44 out45 out46 out47 control	control^	MUX-Array-16-no-INV	wn='wn'	wp='wp'	le='le'
x4	in48-1 in49-1 in50-1 in51-1 in52-1 in53-1 in54-1 in55-1 in56-1 in57-1 in58-1 in59-1 in60-1 in61-1 in62-1 in63-1 in48-2 in49-2 in50-2 in51-2 in52-2 in53-2 in54-2 in55-2 in56-2 in57-2 in58-2 in59-2 in60-2 in61-2 in62-2 in63-2 out48 out49 out50 out51 out52 out53 out54 out55 out56 out57 out58 out59 out60 out61 out62 out63 control	control^	MUX-Array-16-no-INV	wn='wn'	wp='wp'	le='le'
x5	in64-1 in65-1 in66-1 in67-1 in68-1 in69-1 in70-1 in71-1 in72-1 in73-1 in74-1 in75-1 in76-1 in77-1 in78-1 in79-1 in64-2 in65-2 in66-2 in67-2 in68-2 in69-2 in70-2 in71-2 in72-2 in73-2 in74-2 in75-2 in76-2 in77-2 in78-2 in79-2 out64 out65 out66 out67 out68 out69 out70 out71 out72 out73 out74 out75 out76 out77 out78 out79 control	control^	MUX-Array-16-no-INV	wn='wn'	wp='wp'	le='le'
x6	in80-1 in81-1 in82-1 in83-1 in84-1 in85-1 in86-1 in87-1 in88-1 in89-1 in90-1 in91-1 in92-1 in93-1 in94-1 in95-1 in80-2 in81-2 in82-2 in83-2 in84-2 in85-2 in86-2 in87-2 in88-2 in89-2 in90-2 in91-2 in92-2 in93-2 in94-2 in95-2 out80 out81 out82 out83 out84 out85 out86 out87 out88 out89 out90 out91 out92 out93 out94 out95 control	control^	MUX-Array-16-no-INV	wn='wn'	wp='wp'	le='le'
x7	in96-1 in97-1 in98-1 in99-1 in100-1 in101-1 in102-1 in103-1 in104-1 in105-1 in106-1 in107-1 in108-1 in109-1 in110-1 in111-1 in96-2 in97-2 in98-2 in99-2 in100-2 in101-2 in102-2 in103-2 in104-2 in105-2 in106-2 in107-2 in108-2 in109-2 in110-2 in111-2 out96 out97 out98 out99 out100 out101 out102 out103 out104 out105 out106 out107 out108 out109 out110 out111 control	control^	MUX-Array-16-no-INV	wn='wn'	wp='wp'	le='le'
x8	in112-1 in113-1 in114-1 in115-1 in116-1 in117-1 in118-1 in119-1 in120-1 in121-1 in122-1 in123-1 in124-1 in125-1 in126-1 in127-1 in112-2 in113-2 in114-2 in115-2 in116-2 in117-2 in118-2 in119-2 in120-2 in121-2 in122-2 in123-2 in124-2 in125-2 in126-2 in127-2 out112 out113 out114 out115 out116 out117 out118 out119 out120 out121 out122 out123 out124 out125 out126 out127 control	control^	MUX-Array-16-no-INV	wn='wn'	wp='wp'	le='le'
.ends

***Array of 16 inverter-less multiplexers***
.subckt	MUX-Array-16-no-INV	in1-1	in1-2	in1-3	in1-4	in1-5	in1-6	in1-7	in1-8	in1-9	in1-10	in1-11	in1-12	in1-13	in1-14	in1-15	in1-16	in2-1	in2-2	in2-3	in2-4	in2-5	in2-6	in2-7	in2-8	in2-9	in2-10	in2-11	in2-12	in2-13	in2-14	in2-15	in2-16	out1	out2	out3	out4	out5	out6	out7	out8	out9	out10	out11	out12	out13	out14	out15	out16	control	control^	wn=1u	wp=3u	le=0.18u
x1	in1-1	in1-2	in1-3	in1-4	in2-1	in2-2	in2-3	in2-4	out1	out2	out3	out4	control	control^	MUX-Array-4-no-INV	wn='wn'	wp='wp'	le='le'
x2	in1-5	in1-6	in1-7	in1-8	in2-5	in2-6	in2-7	in2-8	out5	out6	out7	out8	control	control^	MUX-Array-4-no-INV	wn='wn'	wp='wp'	le='le'
x3	in1-9	in1-10	in1-11	in1-12	in2-9	in2-10	in2-11	in2-12	out9	out10	out11	out12	control	control^	MUX-Array-4-no-INV	wn='wn'	wp='wp'	le='le'
x4	in1-13	in1-14	in1-15	in1-16	in2-13	in2-14	in2-15	in2-16	out13	out14	out15	out16	control	control^	MUX-Array-4-no-INV	wn='wn'	wp='wp'	le='le'
.ends

***Array of 4 inverter-less multiplexers***
.subckt	MUX-Array-4-no-INV	in1-1	in1-2	in1-3	in1-4	in2-1	in2-2	in2-3	in2-4	out1	out2	out3	out4	control	control^	wn=1u	wp=3u	le=0.18u
x1	in1-1	in2-1	out1	control	control^	MUX-no-INV	wn='wn'	wp='wp'	le='le'
x2	in1-2	in2-2	out2	control	control^	MUX-no-INV	wn='wn'	wp='wp'	le='le'
x3	in1-3	in2-3	out3	control	control^	MUX-no-INV	wn='wn'	wp='wp'	le='le'
x4	in1-4	in2-4	out4	control	control^	MUX-no-INV	wn='wn'	wp='wp'	le='le'
.ends

***20-Transistor Multiplexer without Inverter***
.subckt	MUX-no-INV	in1	in2	out	control	control^	wn=1u	wp=3u	le=0.18u
x1	in1	out	control	control^	TG-m20	wn='wn'	wp='wp'	le='le'
x2	in2	out	control^	control	TG-m20	wn='wn'	wp='wp'	le='le'
.ends

***20-Transistor Transmission Gate***
.subckt	TG-m20	in	out	control	control^	wn=1u	wp=3u	le=0.18u
m1	in	control^	out	vdd	mp18	w=wp	l=le	m=20
m2	out	control	in	0	mn18	w=wn	l=le	m=20
.ends

***20-Transistor Multiplexer***
.subckt	MUX-m20	in1	in2	out	control	wn=1u	wp=3u	le=0.18u
x1	in1	out	control	control^	TG-m20	wn='wn'	wp='wp'	le='le'
x2	in2	out	control^	control	TG-m20	wn='wn'	wp='wp'	le='le'
x3	control	control^	INV-m20	wn='wn'	wp='wp'	le='le'
.ends

***10-Transistor Multiplexer***
.subckt	MUX-m10	in1	in2	out	control	wn=1u	wp=3u	le=0.18u
x1	in1	out	control	control^	TG-m10	wn='wn'	wp='wp'	le='le'
x2	in2	out	control^	control	TG-m10	wn='wn'	wp='wp'	le='le'
x3	control	control^	INV-m10	wn='wn'	wp='wp'	le='le'
.ends

***10-Transistor Transmission Gate***
.subckt	TG-m10	in	out	control	control^	wn=1u	wp=3u	le=0.18u
m1	in	control^	out	vdd	mp18	w=wp	l=le	m=10
m2	out	control	in	0	mn18	w=wn	l=le	m=10
.ends

***10-Transistor Inverter
.subckt	INV-m10	in	out	wn=1u	wp=3u	le=0.18u
m1	out	in	vdd	vdd	mp18	w=wp	l=le	m=10
m2	out	in	0	0	mn18	w=wn	l=le	m=10
.ends

***20-Transistor 2-Input OR***
.subckt	OR2-m20	in1	in2	out	out^	wn=1u	wp=3u	le=0.18u
x1	in1	in2	out^	NOR2-m20	wn='wn'	wp='wp'	le='le'
x2	out^	out	INV-m20	wn='wn'	wp='wp'	le='le'
.ends

***20-Transistor 2-Input NOR***
.subckt	NOR2-m20	in1	in2	out	wn=1u	wp=3u	le=0.18u
m1	a	in2	vdd	vdd	mp18	w='2*wp'	l=le	m=20
m2	out	in1	a	vdd	mp18	w='2*wp'	l=le	m=20
m3	out	in1	0	0	mn18	w=wn	l=le	m=20
m4	out	in2	0	0	mn18	w=wn	l=le	m=20
.ends

***20-Transistor Inverter
.subckt	INV-m20	in	out	wn=1u	wp=3u	le=0.18u
m1	out	in	vdd	vdd	mp18	w=wp	l=le	m=20
m2	out	in	0	0	mn18	w=wn	l=le	m=20
.ends

***10-Transistor 2-Input OR***
.subckt	OR2-m10	in1	in2	out	out^	wn=1u	wp=3u	le=0.18u
x1	in1	in2	out^	NOR2-m10	wn='wn'	wp='wp'	le='le'
x2	out^	out	INV-m10	wn='wn'	wp='wp'	le='le'
.ends

***10-Transistor 2-Input NOR***
.subckt	NOR2-m10	in1	in2	out	wn=1u	wp=3u	le=0.18u
m1	a	in2	vdd	vdd	mp18	w='2*wp'	l=le	m=10
m2	out	in1	a	vdd	mp18	w='2*wp'	l=le	m=10
m3	out	in1	0	0	mn18	w=wn	l=le	m=10
m4	out	in2	0	0	mn18	w=wn	l=le	m=10
.ends

***10-Transistor 2-Input AND***
.subckt	AND2-m10	in1	in2	out	out^	wn=1u	wp=3u	le=0.18u
x1	in1	in2	out^	NAND2-m10	wn='wn'	wp='wp'	le='le'
x2	out^	out	INV-m10	wn='wn'	wp='wp'	le='le'
.ends

***10-Transistor 2-Input NAND***
.subckt	NAND2-m10	in1	in2	out	wn=1u	wp=3u	le=0.18u
m1	out	in1	vdd	vdd	mp18	w=wp	l=le	m=10
m2	out	in2	vdd	vdd	mp18	w=wp	l=le	m=10
m3	out	in1	a	0	mn18	w='2*wn'	l=le	m=10
m4	a	in2	0	0	mn18	w='2*wn'	l=le	m=10
.ends

***20-Transistor 2-Input AND***
.subckt	AND2-m20	in1	in2	out	out^	wn=1u	wp=3u	le=0.18u
x1	in1	in2	out^	NAND2-m20	wn='wn'	wp='wp'	le='le'
x2	out^	out	INV-m20	wn='wn'	wp='wp'	le='le'
.ends

***20-Transistor 2-Input NAND***
.subckt	NAND2-m20	in1	in2	out	wn=1u	wp=3u	le=0.18u
m1	out	in1	vdd	vdd	mp18	w=wp	l=le	m=20
m2	out	in2	vdd	vdd	mp18	w=wp	l=le	m=20
m3	out	in1	a	0	mn18	w='2*wn'	l=le	m=20
m4	a	in2	0	0	mn18	w='2*wn'	l=le	m=20
.ends

***20-Transistor 8-Input AND***
.subckt	AND8-m20	in1	in2	in3	in4	in5	in6	in7	in8	out	out^	wn=1u	wp=3u	le=0.18u
x1	in1	in2	in3	in4	in5	in6	in7	in8	out^	NAND8-m20	wn='wn'	wp='wp'	le='le'
x2	out^	out	INV-m20	wn='wn'	wp='wp'	le='le'
.ends

***20-Transistor 8-Input NAND***
.subckt NAND8-m20	in1	in2	in3	in4	in5	in6	in7	in8	out	wn=1u	wp=3u	le=0.18u
m1	out	in1	vdd	vdd	mp18	w=wp	l=le	m=20
m2	out	in2	vdd	vdd	mp18	w=wp	l=le	m=20
m3	out	in3	vdd	vdd	mp18	w=wp	l=le	m=20
m4	out	in4	vdd	vdd	mp18	w=wp	l=le	m=20
m5	out	in5	vdd	vdd	mp18	w=wp	l=le	m=20
m6	out	in6	vdd	vdd	mp18	w=wp	l=le	m=20
m7	out	in7	vdd	vdd	mp18	w=wp	l=le	m=20
m8	out	in8	vdd	vdd	mp18	w=wp	l=le	m=20

m9	out	in1	a	0	mn18	w='8*wn'	l=le	m=20
m10	a	in2	b	0	mn18	w='8*wn'	l=le	m=20
m11	b	in3	c	0	mn18	w='8*wn'	l=le	m=20
m12	c	in4	d	0	mn18	w='8*wn'	l=le	m=20
m13	d	in5	e	0	mn18	w='8*wn'	l=le	m=20
m14	e	in6	f	0	mn18	w='8*wn'	l=le	m=20
m15	f	in7	g	0	mn18	w='8*wn'	l=le	m=20
m16	g	in8	0	0	mn18	w='8*wn'	l=le	m=20
.ends

******Include
.include	'./GAP.inc'
*.include	'./RAM.inc'

.end
